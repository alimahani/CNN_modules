module bc_pe(
  input         clock,
  input         reset,
  input  [15:0] io_ho_input,
  input  [31:0] io_ve_input,
  input         io_input_valid,
  input         io_iormac,
  output [31:0] io_ve_out,
  output [15:0] io_ho_out,
  output [31:0] io_res_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mac; // @[bc_pe.scala 30:23]
  reg [15:0] ho_reg; // @[bc_pe.scala 31:23]
  reg [31:0] ve_reg; // @[bc_pe.scala 32:23]
  reg  REG; // @[bc_pe.scala 37:42]
  wire  _T_1 = io_input_valid & ~REG; // @[bc_pe.scala 37:31]
  wire [47:0] _mac_T = io_ho_input * io_ve_input; // @[bc_pe.scala 44:39]
  wire [47:0] _GEN_3 = {{16'd0}, mac}; // @[bc_pe.scala 44:24]
  wire [47:0] _mac_T_2 = _GEN_3 + _mac_T; // @[bc_pe.scala 44:24]
  wire [47:0] _GEN_0 = _T_1 ? _mac_T_2 : {{16'd0}, mac}; // @[bc_pe.scala 42:46 44:17 30:23]
  wire [47:0] _GEN_4 = reset ? 48'h0 : _GEN_0; // @[bc_pe.scala 30:{23,23}]
  assign io_ve_out = io_iormac ? ve_reg : mac; // @[bc_pe.scala 51:20]
  assign io_ho_out = ho_reg; // @[bc_pe.scala 52:14]
  assign io_res_out = mac; // @[bc_pe.scala 50:14]
  always @(posedge clock) begin
    mac <= _GEN_4[31:0]; // @[bc_pe.scala 30:{23,23}]
    if (reset) begin // @[bc_pe.scala 31:23]
      ho_reg <= 16'h0; // @[bc_pe.scala 31:23]
    end else if (_T_1) begin // @[bc_pe.scala 42:46]
      ho_reg <= io_ho_input; // @[bc_pe.scala 45:17]
    end
    if (reset) begin // @[bc_pe.scala 32:23]
      ve_reg <= 32'h0; // @[bc_pe.scala 32:23]
    end else if (_T_1) begin // @[bc_pe.scala 42:46]
      ve_reg <= io_ve_input; // @[bc_pe.scala 46:17]
    end
    REG <= io_input_valid; // @[bc_pe.scala 37:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mac = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ho_reg = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  ve_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  REG = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module bc_mmul(
  input         clock,
  input         reset,
  input  [15:0] io_x_input_0,
  input  [15:0] io_x_input_1,
  input  [15:0] io_x_input_2,
  input  [15:0] io_x_input_3,
  input  [15:0] io_x_input_4,
  input  [15:0] io_x_input_5,
  input  [15:0] io_x_input_6,
  input  [15:0] io_x_input_7,
  input  [15:0] io_x_input_8,
  input  [15:0] io_x_input_9,
  input  [15:0] io_x_input_10,
  input  [15:0] io_x_input_11,
  input  [15:0] io_x_input_12,
  input  [15:0] io_x_input_13,
  input  [15:0] io_x_input_14,
  input  [15:0] io_x_input_15,
  input  [15:0] io_x_input_16,
  input  [15:0] io_x_input_17,
  input  [15:0] io_x_input_18,
  input  [15:0] io_x_input_19,
  input  [15:0] io_x_input_20,
  input  [15:0] io_x_input_21,
  input  [15:0] io_x_input_22,
  input  [15:0] io_x_input_23,
  input  [15:0] io_x_input_24,
  input  [15:0] io_x_input_25,
  input  [15:0] io_x_input_26,
  input  [15:0] io_x_input_27,
  input  [15:0] io_x_input_28,
  input  [15:0] io_x_input_29,
  input  [15:0] io_x_input_30,
  input  [15:0] io_x_input_31,
  input  [31:0] io_w_input_0,
  input  [31:0] io_w_input_1,
  input  [31:0] io_w_input_2,
  input  [31:0] io_w_input_3,
  input  [31:0] io_w_input_4,
  input  [31:0] io_w_input_5,
  input  [31:0] io_w_input_6,
  input  [31:0] io_w_input_7,
  input  [31:0] io_w_input_8,
  input  [31:0] io_w_input_9,
  input  [31:0] io_w_input_10,
  input  [31:0] io_w_input_11,
  input  [31:0] io_w_input_12,
  input  [31:0] io_w_input_13,
  input  [31:0] io_w_input_14,
  input  [31:0] io_w_input_15,
  input  [31:0] io_w_input_16,
  input  [31:0] io_w_input_17,
  input  [31:0] io_w_input_18,
  input  [31:0] io_w_input_19,
  input  [31:0] io_w_input_20,
  input  [31:0] io_w_input_21,
  input  [31:0] io_w_input_22,
  input  [31:0] io_w_input_23,
  input  [31:0] io_w_input_24,
  input  [31:0] io_w_input_25,
  input  [31:0] io_w_input_26,
  input  [31:0] io_w_input_27,
  input  [31:0] io_w_input_28,
  input  [31:0] io_w_input_29,
  input  [31:0] io_w_input_30,
  input  [31:0] io_w_input_31,
  input         io_input_valid_0,
  input         io_input_valid_1,
  input         io_input_valid_2,
  input         io_input_valid_3,
  input         io_input_valid_4,
  input         io_input_valid_5,
  input         io_input_valid_6,
  input         io_input_valid_7,
  input         io_input_valid_8,
  input         io_input_valid_9,
  input         io_input_valid_10,
  input         io_input_valid_11,
  input         io_input_valid_12,
  input         io_input_valid_13,
  input         io_input_valid_14,
  input         io_input_valid_15,
  input         io_input_valid_16,
  input         io_input_valid_17,
  input         io_input_valid_18,
  input         io_input_valid_19,
  input         io_input_valid_20,
  input         io_input_valid_21,
  input         io_input_valid_22,
  input         io_input_valid_23,
  input         io_input_valid_24,
  input         io_input_valid_25,
  input         io_input_valid_26,
  input         io_input_valid_27,
  input         io_input_valid_28,
  input         io_input_valid_29,
  input         io_input_valid_30,
  input         io_input_valid_31,
  input         io_input_valid_32,
  input         io_input_valid_33,
  input         io_input_valid_34,
  input         io_input_valid_35,
  input         io_input_valid_36,
  input         io_input_valid_37,
  input         io_input_valid_38,
  input         io_input_valid_39,
  input         io_input_valid_40,
  input         io_input_valid_41,
  input         io_input_valid_42,
  input         io_input_valid_43,
  input         io_input_valid_44,
  input         io_input_valid_45,
  input         io_input_valid_46,
  input         io_input_valid_47,
  input         io_input_valid_48,
  input         io_input_valid_49,
  input         io_input_valid_50,
  input         io_input_valid_51,
  input         io_input_valid_52,
  input         io_input_valid_53,
  input         io_input_valid_54,
  input         io_input_valid_55,
  input         io_input_valid_56,
  input         io_input_valid_57,
  input         io_input_valid_58,
  input         io_input_valid_59,
  input         io_input_valid_60,
  input         io_input_valid_61,
  input         io_input_valid_62,
  input         io_input_valid_63,
  input         io_input_valid_64,
  input         io_input_valid_65,
  input         io_input_valid_66,
  input         io_input_valid_67,
  input         io_input_valid_68,
  input         io_input_valid_69,
  input         io_input_valid_70,
  input         io_input_valid_71,
  input         io_input_valid_72,
  input         io_input_valid_73,
  input         io_input_valid_74,
  input         io_input_valid_75,
  input         io_input_valid_76,
  input         io_input_valid_77,
  input         io_input_valid_78,
  input         io_input_valid_79,
  input         io_input_valid_80,
  input         io_input_valid_81,
  input         io_input_valid_82,
  input         io_input_valid_83,
  input         io_input_valid_84,
  input         io_input_valid_85,
  input         io_input_valid_86,
  input         io_input_valid_87,
  input         io_input_valid_88,
  input         io_input_valid_89,
  input         io_input_valid_90,
  input         io_input_valid_91,
  input         io_input_valid_92,
  input         io_input_valid_93,
  input         io_input_valid_94,
  input         io_input_valid_95,
  input         io_input_valid_96,
  input         io_input_valid_97,
  input         io_input_valid_98,
  input         io_input_valid_99,
  input         io_input_valid_100,
  input         io_input_valid_101,
  input         io_input_valid_102,
  input         io_input_valid_103,
  input         io_input_valid_104,
  input         io_input_valid_105,
  input         io_input_valid_106,
  input         io_input_valid_107,
  input         io_input_valid_108,
  input         io_input_valid_109,
  input         io_input_valid_110,
  input         io_input_valid_111,
  input         io_input_valid_112,
  input         io_input_valid_113,
  input         io_input_valid_114,
  input         io_input_valid_115,
  input         io_input_valid_116,
  input         io_input_valid_117,
  input         io_input_valid_118,
  input         io_input_valid_119,
  input         io_input_valid_120,
  input         io_input_valid_121,
  input         io_input_valid_122,
  input         io_input_valid_123,
  input         io_input_valid_124,
  input         io_input_valid_125,
  input         io_input_valid_126,
  input         io_input_valid_127,
  input         io_input_valid_128,
  input         io_input_valid_129,
  input         io_input_valid_130,
  input         io_input_valid_131,
  input         io_input_valid_132,
  input         io_input_valid_133,
  input         io_input_valid_134,
  input         io_input_valid_135,
  input         io_input_valid_136,
  input         io_input_valid_137,
  input         io_input_valid_138,
  input         io_input_valid_139,
  input         io_input_valid_140,
  input         io_input_valid_141,
  input         io_input_valid_142,
  input         io_input_valid_143,
  input         io_input_valid_144,
  input         io_input_valid_145,
  input         io_input_valid_146,
  input         io_input_valid_147,
  input         io_input_valid_148,
  input         io_input_valid_149,
  input         io_input_valid_150,
  input         io_input_valid_151,
  input         io_input_valid_152,
  input         io_input_valid_153,
  input         io_input_valid_154,
  input         io_input_valid_155,
  input         io_input_valid_156,
  input         io_input_valid_157,
  input         io_input_valid_158,
  input         io_input_valid_159,
  input         io_input_valid_160,
  input         io_input_valid_161,
  input         io_input_valid_162,
  input         io_input_valid_163,
  input         io_input_valid_164,
  input         io_input_valid_165,
  input         io_input_valid_166,
  input         io_input_valid_167,
  input         io_input_valid_168,
  input         io_input_valid_169,
  input         io_input_valid_170,
  input         io_input_valid_171,
  input         io_input_valid_172,
  input         io_input_valid_173,
  input         io_input_valid_174,
  input         io_input_valid_175,
  input         io_input_valid_176,
  input         io_input_valid_177,
  input         io_input_valid_178,
  input         io_input_valid_179,
  input         io_input_valid_180,
  input         io_input_valid_181,
  input         io_input_valid_182,
  input         io_input_valid_183,
  input         io_input_valid_184,
  input         io_input_valid_185,
  input         io_input_valid_186,
  input         io_input_valid_187,
  input         io_input_valid_188,
  input         io_input_valid_189,
  input         io_input_valid_190,
  input         io_input_valid_191,
  input         io_input_valid_192,
  input         io_input_valid_193,
  input         io_input_valid_194,
  input         io_input_valid_195,
  input         io_input_valid_196,
  input         io_input_valid_197,
  input         io_input_valid_198,
  input         io_input_valid_199,
  input         io_input_valid_200,
  input         io_input_valid_201,
  input         io_input_valid_202,
  input         io_input_valid_203,
  input         io_input_valid_204,
  input         io_input_valid_205,
  input         io_input_valid_206,
  input         io_input_valid_207,
  input         io_input_valid_208,
  input         io_input_valid_209,
  input         io_input_valid_210,
  input         io_input_valid_211,
  input         io_input_valid_212,
  input         io_input_valid_213,
  input         io_input_valid_214,
  input         io_input_valid_215,
  input         io_input_valid_216,
  input         io_input_valid_217,
  input         io_input_valid_218,
  input         io_input_valid_219,
  input         io_input_valid_220,
  input         io_input_valid_221,
  input         io_input_valid_222,
  input         io_input_valid_223,
  input         io_input_valid_224,
  input         io_input_valid_225,
  input         io_input_valid_226,
  input         io_input_valid_227,
  input         io_input_valid_228,
  input         io_input_valid_229,
  input         io_input_valid_230,
  input         io_input_valid_231,
  input         io_input_valid_232,
  input         io_input_valid_233,
  input         io_input_valid_234,
  input         io_input_valid_235,
  input         io_input_valid_236,
  input         io_input_valid_237,
  input         io_input_valid_238,
  input         io_input_valid_239,
  input         io_input_valid_240,
  input         io_input_valid_241,
  input         io_input_valid_242,
  input         io_input_valid_243,
  input         io_input_valid_244,
  input         io_input_valid_245,
  input         io_input_valid_246,
  input         io_input_valid_247,
  input         io_input_valid_248,
  input         io_input_valid_249,
  input         io_input_valid_250,
  input         io_input_valid_251,
  input         io_input_valid_252,
  input         io_input_valid_253,
  input         io_input_valid_254,
  input         io_input_valid_255,
  input         io_input_valid_256,
  input         io_input_valid_257,
  input         io_input_valid_258,
  input         io_input_valid_259,
  input         io_input_valid_260,
  input         io_input_valid_261,
  input         io_input_valid_262,
  input         io_input_valid_263,
  input         io_input_valid_264,
  input         io_input_valid_265,
  input         io_input_valid_266,
  input         io_input_valid_267,
  input         io_input_valid_268,
  input         io_input_valid_269,
  input         io_input_valid_270,
  input         io_input_valid_271,
  input         io_input_valid_272,
  input         io_input_valid_273,
  input         io_input_valid_274,
  input         io_input_valid_275,
  input         io_input_valid_276,
  input         io_input_valid_277,
  input         io_input_valid_278,
  input         io_input_valid_279,
  input         io_input_valid_280,
  input         io_input_valid_281,
  input         io_input_valid_282,
  input         io_input_valid_283,
  input         io_input_valid_284,
  input         io_input_valid_285,
  input         io_input_valid_286,
  input         io_input_valid_287,
  input         io_input_valid_288,
  input         io_input_valid_289,
  input         io_input_valid_290,
  input         io_input_valid_291,
  input         io_input_valid_292,
  input         io_input_valid_293,
  input         io_input_valid_294,
  input         io_input_valid_295,
  input         io_input_valid_296,
  input         io_input_valid_297,
  input         io_input_valid_298,
  input         io_input_valid_299,
  input         io_input_valid_300,
  input         io_input_valid_301,
  input         io_input_valid_302,
  input         io_input_valid_303,
  input         io_input_valid_304,
  input         io_input_valid_305,
  input         io_input_valid_306,
  input         io_input_valid_307,
  input         io_input_valid_308,
  input         io_input_valid_309,
  input         io_input_valid_310,
  input         io_input_valid_311,
  input         io_input_valid_312,
  input         io_input_valid_313,
  input         io_input_valid_314,
  input         io_input_valid_315,
  input         io_input_valid_316,
  input         io_input_valid_317,
  input         io_input_valid_318,
  input         io_input_valid_319,
  input         io_input_valid_320,
  input         io_input_valid_321,
  input         io_input_valid_322,
  input         io_input_valid_323,
  input         io_input_valid_324,
  input         io_input_valid_325,
  input         io_input_valid_326,
  input         io_input_valid_327,
  input         io_input_valid_328,
  input         io_input_valid_329,
  input         io_input_valid_330,
  input         io_input_valid_331,
  input         io_input_valid_332,
  input         io_input_valid_333,
  input         io_input_valid_334,
  input         io_input_valid_335,
  input         io_input_valid_336,
  input         io_input_valid_337,
  input         io_input_valid_338,
  input         io_input_valid_339,
  input         io_input_valid_340,
  input         io_input_valid_341,
  input         io_input_valid_342,
  input         io_input_valid_343,
  input         io_input_valid_344,
  input         io_input_valid_345,
  input         io_input_valid_346,
  input         io_input_valid_347,
  input         io_input_valid_348,
  input         io_input_valid_349,
  input         io_input_valid_350,
  input         io_input_valid_351,
  input         io_input_valid_352,
  input         io_input_valid_353,
  input         io_input_valid_354,
  input         io_input_valid_355,
  input         io_input_valid_356,
  input         io_input_valid_357,
  input         io_input_valid_358,
  input         io_input_valid_359,
  input         io_input_valid_360,
  input         io_input_valid_361,
  input         io_input_valid_362,
  input         io_input_valid_363,
  input         io_input_valid_364,
  input         io_input_valid_365,
  input         io_input_valid_366,
  input         io_input_valid_367,
  input         io_input_valid_368,
  input         io_input_valid_369,
  input         io_input_valid_370,
  input         io_input_valid_371,
  input         io_input_valid_372,
  input         io_input_valid_373,
  input         io_input_valid_374,
  input         io_input_valid_375,
  input         io_input_valid_376,
  input         io_input_valid_377,
  input         io_input_valid_378,
  input         io_input_valid_379,
  input         io_input_valid_380,
  input         io_input_valid_381,
  input         io_input_valid_382,
  input         io_input_valid_383,
  input         io_input_valid_384,
  input         io_input_valid_385,
  input         io_input_valid_386,
  input         io_input_valid_387,
  input         io_input_valid_388,
  input         io_input_valid_389,
  input         io_input_valid_390,
  input         io_input_valid_391,
  input         io_input_valid_392,
  input         io_input_valid_393,
  input         io_input_valid_394,
  input         io_input_valid_395,
  input         io_input_valid_396,
  input         io_input_valid_397,
  input         io_input_valid_398,
  input         io_input_valid_399,
  input         io_input_valid_400,
  input         io_input_valid_401,
  input         io_input_valid_402,
  input         io_input_valid_403,
  input         io_input_valid_404,
  input         io_input_valid_405,
  input         io_input_valid_406,
  input         io_input_valid_407,
  input         io_input_valid_408,
  input         io_input_valid_409,
  input         io_input_valid_410,
  input         io_input_valid_411,
  input         io_input_valid_412,
  input         io_input_valid_413,
  input         io_input_valid_414,
  input         io_input_valid_415,
  input         io_input_valid_416,
  input         io_input_valid_417,
  input         io_input_valid_418,
  input         io_input_valid_419,
  input         io_input_valid_420,
  input         io_input_valid_421,
  input         io_input_valid_422,
  input         io_input_valid_423,
  input         io_input_valid_424,
  input         io_input_valid_425,
  input         io_input_valid_426,
  input         io_input_valid_427,
  input         io_input_valid_428,
  input         io_input_valid_429,
  input         io_input_valid_430,
  input         io_input_valid_431,
  input         io_input_valid_432,
  input         io_input_valid_433,
  input         io_input_valid_434,
  input         io_input_valid_435,
  input         io_input_valid_436,
  input         io_input_valid_437,
  input         io_input_valid_438,
  input         io_input_valid_439,
  input         io_input_valid_440,
  input         io_input_valid_441,
  input         io_input_valid_442,
  input         io_input_valid_443,
  input         io_input_valid_444,
  input         io_input_valid_445,
  input         io_input_valid_446,
  input         io_input_valid_447,
  input         io_input_valid_448,
  input         io_input_valid_449,
  input         io_input_valid_450,
  input         io_input_valid_451,
  input         io_input_valid_452,
  input         io_input_valid_453,
  input         io_input_valid_454,
  input         io_input_valid_455,
  input         io_input_valid_456,
  input         io_input_valid_457,
  input         io_input_valid_458,
  input         io_input_valid_459,
  input         io_input_valid_460,
  input         io_input_valid_461,
  input         io_input_valid_462,
  input         io_input_valid_463,
  input         io_input_valid_464,
  input         io_input_valid_465,
  input         io_input_valid_466,
  input         io_input_valid_467,
  input         io_input_valid_468,
  input         io_input_valid_469,
  input         io_input_valid_470,
  input         io_input_valid_471,
  input         io_input_valid_472,
  input         io_input_valid_473,
  input         io_input_valid_474,
  input         io_input_valid_475,
  input         io_input_valid_476,
  input         io_input_valid_477,
  input         io_input_valid_478,
  input         io_input_valid_479,
  input         io_input_valid_480,
  input         io_input_valid_481,
  input         io_input_valid_482,
  input         io_input_valid_483,
  input         io_input_valid_484,
  input         io_input_valid_485,
  input         io_input_valid_486,
  input         io_input_valid_487,
  input         io_input_valid_488,
  input         io_input_valid_489,
  input         io_input_valid_490,
  input         io_input_valid_491,
  input         io_input_valid_492,
  input         io_input_valid_493,
  input         io_input_valid_494,
  input         io_input_valid_495,
  input         io_input_valid_496,
  input         io_input_valid_497,
  input         io_input_valid_498,
  input         io_input_valid_499,
  input         io_input_valid_500,
  input         io_input_valid_501,
  input         io_input_valid_502,
  input         io_input_valid_503,
  input         io_input_valid_504,
  input         io_input_valid_505,
  input         io_input_valid_506,
  input         io_input_valid_507,
  input         io_input_valid_508,
  input         io_input_valid_509,
  input         io_input_valid_510,
  input         io_input_valid_511,
  input         io_input_valid_512,
  input         io_input_valid_513,
  input         io_input_valid_514,
  input         io_input_valid_515,
  input         io_input_valid_516,
  input         io_input_valid_517,
  input         io_input_valid_518,
  input         io_input_valid_519,
  input         io_input_valid_520,
  input         io_input_valid_521,
  input         io_input_valid_522,
  input         io_input_valid_523,
  input         io_input_valid_524,
  input         io_input_valid_525,
  input         io_input_valid_526,
  input         io_input_valid_527,
  input         io_input_valid_528,
  input         io_input_valid_529,
  input         io_input_valid_530,
  input         io_input_valid_531,
  input         io_input_valid_532,
  input         io_input_valid_533,
  input         io_input_valid_534,
  input         io_input_valid_535,
  input         io_input_valid_536,
  input         io_input_valid_537,
  input         io_input_valid_538,
  input         io_input_valid_539,
  input         io_input_valid_540,
  input         io_input_valid_541,
  input         io_input_valid_542,
  input         io_input_valid_543,
  input         io_input_valid_544,
  input         io_input_valid_545,
  input         io_input_valid_546,
  input         io_input_valid_547,
  input         io_input_valid_548,
  input         io_input_valid_549,
  input         io_input_valid_550,
  input         io_input_valid_551,
  input         io_input_valid_552,
  input         io_input_valid_553,
  input         io_input_valid_554,
  input         io_input_valid_555,
  input         io_input_valid_556,
  input         io_input_valid_557,
  input         io_input_valid_558,
  input         io_input_valid_559,
  input         io_input_valid_560,
  input         io_input_valid_561,
  input         io_input_valid_562,
  input         io_input_valid_563,
  input         io_input_valid_564,
  input         io_input_valid_565,
  input         io_input_valid_566,
  input         io_input_valid_567,
  input         io_input_valid_568,
  input         io_input_valid_569,
  input         io_input_valid_570,
  input         io_input_valid_571,
  input         io_input_valid_572,
  input         io_input_valid_573,
  input         io_input_valid_574,
  input         io_input_valid_575,
  input         io_input_valid_576,
  input         io_input_valid_577,
  input         io_input_valid_578,
  input         io_input_valid_579,
  input         io_input_valid_580,
  input         io_input_valid_581,
  input         io_input_valid_582,
  input         io_input_valid_583,
  input         io_input_valid_584,
  input         io_input_valid_585,
  input         io_input_valid_586,
  input         io_input_valid_587,
  input         io_input_valid_588,
  input         io_input_valid_589,
  input         io_input_valid_590,
  input         io_input_valid_591,
  input         io_input_valid_592,
  input         io_input_valid_593,
  input         io_input_valid_594,
  input         io_input_valid_595,
  input         io_input_valid_596,
  input         io_input_valid_597,
  input         io_input_valid_598,
  input         io_input_valid_599,
  input         io_input_valid_600,
  input         io_input_valid_601,
  input         io_input_valid_602,
  input         io_input_valid_603,
  input         io_input_valid_604,
  input         io_input_valid_605,
  input         io_input_valid_606,
  input         io_input_valid_607,
  input         io_input_valid_608,
  input         io_input_valid_609,
  input         io_input_valid_610,
  input         io_input_valid_611,
  input         io_input_valid_612,
  input         io_input_valid_613,
  input         io_input_valid_614,
  input         io_input_valid_615,
  input         io_input_valid_616,
  input         io_input_valid_617,
  input         io_input_valid_618,
  input         io_input_valid_619,
  input         io_input_valid_620,
  input         io_input_valid_621,
  input         io_input_valid_622,
  input         io_input_valid_623,
  input         io_input_valid_624,
  input         io_input_valid_625,
  input         io_input_valid_626,
  input         io_input_valid_627,
  input         io_input_valid_628,
  input         io_input_valid_629,
  input         io_input_valid_630,
  input         io_input_valid_631,
  input         io_input_valid_632,
  input         io_input_valid_633,
  input         io_input_valid_634,
  input         io_input_valid_635,
  input         io_input_valid_636,
  input         io_input_valid_637,
  input         io_input_valid_638,
  input         io_input_valid_639,
  input         io_input_valid_640,
  input         io_input_valid_641,
  input         io_input_valid_642,
  input         io_input_valid_643,
  input         io_input_valid_644,
  input         io_input_valid_645,
  input         io_input_valid_646,
  input         io_input_valid_647,
  input         io_input_valid_648,
  input         io_input_valid_649,
  input         io_input_valid_650,
  input         io_input_valid_651,
  input         io_input_valid_652,
  input         io_input_valid_653,
  input         io_input_valid_654,
  input         io_input_valid_655,
  input         io_input_valid_656,
  input         io_input_valid_657,
  input         io_input_valid_658,
  input         io_input_valid_659,
  input         io_input_valid_660,
  input         io_input_valid_661,
  input         io_input_valid_662,
  input         io_input_valid_663,
  input         io_input_valid_664,
  input         io_input_valid_665,
  input         io_input_valid_666,
  input         io_input_valid_667,
  input         io_input_valid_668,
  input         io_input_valid_669,
  input         io_input_valid_670,
  input         io_input_valid_671,
  input         io_input_valid_672,
  input         io_input_valid_673,
  input         io_input_valid_674,
  input         io_input_valid_675,
  input         io_input_valid_676,
  input         io_input_valid_677,
  input         io_input_valid_678,
  input         io_input_valid_679,
  input         io_input_valid_680,
  input         io_input_valid_681,
  input         io_input_valid_682,
  input         io_input_valid_683,
  input         io_input_valid_684,
  input         io_input_valid_685,
  input         io_input_valid_686,
  input         io_input_valid_687,
  input         io_input_valid_688,
  input         io_input_valid_689,
  input         io_input_valid_690,
  input         io_input_valid_691,
  input         io_input_valid_692,
  input         io_input_valid_693,
  input         io_input_valid_694,
  input         io_input_valid_695,
  input         io_input_valid_696,
  input         io_input_valid_697,
  input         io_input_valid_698,
  input         io_input_valid_699,
  input         io_input_valid_700,
  input         io_input_valid_701,
  input         io_input_valid_702,
  input         io_input_valid_703,
  input         io_input_valid_704,
  input         io_input_valid_705,
  input         io_input_valid_706,
  input         io_input_valid_707,
  input         io_input_valid_708,
  input         io_input_valid_709,
  input         io_input_valid_710,
  input         io_input_valid_711,
  input         io_input_valid_712,
  input         io_input_valid_713,
  input         io_input_valid_714,
  input         io_input_valid_715,
  input         io_input_valid_716,
  input         io_input_valid_717,
  input         io_input_valid_718,
  input         io_input_valid_719,
  input         io_input_valid_720,
  input         io_input_valid_721,
  input         io_input_valid_722,
  input         io_input_valid_723,
  input         io_input_valid_724,
  input         io_input_valid_725,
  input         io_input_valid_726,
  input         io_input_valid_727,
  input         io_input_valid_728,
  input         io_input_valid_729,
  input         io_input_valid_730,
  input         io_input_valid_731,
  input         io_input_valid_732,
  input         io_input_valid_733,
  input         io_input_valid_734,
  input         io_input_valid_735,
  input         io_input_valid_736,
  input         io_input_valid_737,
  input         io_input_valid_738,
  input         io_input_valid_739,
  input         io_input_valid_740,
  input         io_input_valid_741,
  input         io_input_valid_742,
  input         io_input_valid_743,
  input         io_input_valid_744,
  input         io_input_valid_745,
  input         io_input_valid_746,
  input         io_input_valid_747,
  input         io_input_valid_748,
  input         io_input_valid_749,
  input         io_input_valid_750,
  input         io_input_valid_751,
  input         io_input_valid_752,
  input         io_input_valid_753,
  input         io_input_valid_754,
  input         io_input_valid_755,
  input         io_input_valid_756,
  input         io_input_valid_757,
  input         io_input_valid_758,
  input         io_input_valid_759,
  input         io_input_valid_760,
  input         io_input_valid_761,
  input         io_input_valid_762,
  input         io_input_valid_763,
  input         io_input_valid_764,
  input         io_input_valid_765,
  input         io_input_valid_766,
  input         io_input_valid_767,
  input         io_input_valid_768,
  input         io_input_valid_769,
  input         io_input_valid_770,
  input         io_input_valid_771,
  input         io_input_valid_772,
  input         io_input_valid_773,
  input         io_input_valid_774,
  input         io_input_valid_775,
  input         io_input_valid_776,
  input         io_input_valid_777,
  input         io_input_valid_778,
  input         io_input_valid_779,
  input         io_input_valid_780,
  input         io_input_valid_781,
  input         io_input_valid_782,
  input         io_input_valid_783,
  input         io_input_valid_784,
  input         io_input_valid_785,
  input         io_input_valid_786,
  input         io_input_valid_787,
  input         io_input_valid_788,
  input         io_input_valid_789,
  input         io_input_valid_790,
  input         io_input_valid_791,
  input         io_input_valid_792,
  input         io_input_valid_793,
  input         io_input_valid_794,
  input         io_input_valid_795,
  input         io_input_valid_796,
  input         io_input_valid_797,
  input         io_input_valid_798,
  input         io_input_valid_799,
  input         io_input_valid_800,
  input         io_input_valid_801,
  input         io_input_valid_802,
  input         io_input_valid_803,
  input         io_input_valid_804,
  input         io_input_valid_805,
  input         io_input_valid_806,
  input         io_input_valid_807,
  input         io_input_valid_808,
  input         io_input_valid_809,
  input         io_input_valid_810,
  input         io_input_valid_811,
  input         io_input_valid_812,
  input         io_input_valid_813,
  input         io_input_valid_814,
  input         io_input_valid_815,
  input         io_input_valid_816,
  input         io_input_valid_817,
  input         io_input_valid_818,
  input         io_input_valid_819,
  input         io_input_valid_820,
  input         io_input_valid_821,
  input         io_input_valid_822,
  input         io_input_valid_823,
  input         io_input_valid_824,
  input         io_input_valid_825,
  input         io_input_valid_826,
  input         io_input_valid_827,
  input         io_input_valid_828,
  input         io_input_valid_829,
  input         io_input_valid_830,
  input         io_input_valid_831,
  input         io_input_valid_832,
  input         io_input_valid_833,
  input         io_input_valid_834,
  input         io_input_valid_835,
  input         io_input_valid_836,
  input         io_input_valid_837,
  input         io_input_valid_838,
  input         io_input_valid_839,
  input         io_input_valid_840,
  input         io_input_valid_841,
  input         io_input_valid_842,
  input         io_input_valid_843,
  input         io_input_valid_844,
  input         io_input_valid_845,
  input         io_input_valid_846,
  input         io_input_valid_847,
  input         io_input_valid_848,
  input         io_input_valid_849,
  input         io_input_valid_850,
  input         io_input_valid_851,
  input         io_input_valid_852,
  input         io_input_valid_853,
  input         io_input_valid_854,
  input         io_input_valid_855,
  input         io_input_valid_856,
  input         io_input_valid_857,
  input         io_input_valid_858,
  input         io_input_valid_859,
  input         io_input_valid_860,
  input         io_input_valid_861,
  input         io_input_valid_862,
  input         io_input_valid_863,
  input         io_input_valid_864,
  input         io_input_valid_865,
  input         io_input_valid_866,
  input         io_input_valid_867,
  input         io_input_valid_868,
  input         io_input_valid_869,
  input         io_input_valid_870,
  input         io_input_valid_871,
  input         io_input_valid_872,
  input         io_input_valid_873,
  input         io_input_valid_874,
  input         io_input_valid_875,
  input         io_input_valid_876,
  input         io_input_valid_877,
  input         io_input_valid_878,
  input         io_input_valid_879,
  input         io_input_valid_880,
  input         io_input_valid_881,
  input         io_input_valid_882,
  input         io_input_valid_883,
  input         io_input_valid_884,
  input         io_input_valid_885,
  input         io_input_valid_886,
  input         io_input_valid_887,
  input         io_input_valid_888,
  input         io_input_valid_889,
  input         io_input_valid_890,
  input         io_input_valid_891,
  input         io_input_valid_892,
  input         io_input_valid_893,
  input         io_input_valid_894,
  input         io_input_valid_895,
  input         io_input_valid_896,
  input         io_input_valid_897,
  input         io_input_valid_898,
  input         io_input_valid_899,
  input         io_input_valid_900,
  input         io_input_valid_901,
  input         io_input_valid_902,
  input         io_input_valid_903,
  input         io_input_valid_904,
  input         io_input_valid_905,
  input         io_input_valid_906,
  input         io_input_valid_907,
  input         io_input_valid_908,
  input         io_input_valid_909,
  input         io_input_valid_910,
  input         io_input_valid_911,
  input         io_input_valid_912,
  input         io_input_valid_913,
  input         io_input_valid_914,
  input         io_input_valid_915,
  input         io_input_valid_916,
  input         io_input_valid_917,
  input         io_input_valid_918,
  input         io_input_valid_919,
  input         io_input_valid_920,
  input         io_input_valid_921,
  input         io_input_valid_922,
  input         io_input_valid_923,
  input         io_input_valid_924,
  input         io_input_valid_925,
  input         io_input_valid_926,
  input         io_input_valid_927,
  input         io_input_valid_928,
  input         io_input_valid_929,
  input         io_input_valid_930,
  input         io_input_valid_931,
  input         io_input_valid_932,
  input         io_input_valid_933,
  input         io_input_valid_934,
  input         io_input_valid_935,
  input         io_input_valid_936,
  input         io_input_valid_937,
  input         io_input_valid_938,
  input         io_input_valid_939,
  input         io_input_valid_940,
  input         io_input_valid_941,
  input         io_input_valid_942,
  input         io_input_valid_943,
  input         io_input_valid_944,
  input         io_input_valid_945,
  input         io_input_valid_946,
  input         io_input_valid_947,
  input         io_input_valid_948,
  input         io_input_valid_949,
  input         io_input_valid_950,
  input         io_input_valid_951,
  input         io_input_valid_952,
  input         io_input_valid_953,
  input         io_input_valid_954,
  input         io_input_valid_955,
  input         io_input_valid_956,
  input         io_input_valid_957,
  input         io_input_valid_958,
  input         io_input_valid_959,
  input         io_input_valid_960,
  input         io_input_valid_961,
  input         io_input_valid_962,
  input         io_input_valid_963,
  input         io_input_valid_964,
  input         io_input_valid_965,
  input         io_input_valid_966,
  input         io_input_valid_967,
  input         io_input_valid_968,
  input         io_input_valid_969,
  input         io_input_valid_970,
  input         io_input_valid_971,
  input         io_input_valid_972,
  input         io_input_valid_973,
  input         io_input_valid_974,
  input         io_input_valid_975,
  input         io_input_valid_976,
  input         io_input_valid_977,
  input         io_input_valid_978,
  input         io_input_valid_979,
  input         io_input_valid_980,
  input         io_input_valid_981,
  input         io_input_valid_982,
  input         io_input_valid_983,
  input         io_input_valid_984,
  input         io_input_valid_985,
  input         io_input_valid_986,
  input         io_input_valid_987,
  input         io_input_valid_988,
  input         io_input_valid_989,
  input         io_input_valid_990,
  input         io_input_valid_991,
  input         io_input_valid_992,
  input         io_input_valid_993,
  input         io_input_valid_994,
  input         io_input_valid_995,
  input         io_input_valid_996,
  input         io_input_valid_997,
  input         io_input_valid_998,
  input         io_input_valid_999,
  input         io_input_valid_1000,
  input         io_input_valid_1001,
  input         io_input_valid_1002,
  input         io_input_valid_1003,
  input         io_input_valid_1004,
  input         io_input_valid_1005,
  input         io_input_valid_1006,
  input         io_input_valid_1007,
  input         io_input_valid_1008,
  input         io_input_valid_1009,
  input         io_input_valid_1010,
  input         io_input_valid_1011,
  input         io_input_valid_1012,
  input         io_input_valid_1013,
  input         io_input_valid_1014,
  input         io_input_valid_1015,
  input         io_input_valid_1016,
  input         io_input_valid_1017,
  input         io_input_valid_1018,
  input         io_input_valid_1019,
  input         io_input_valid_1020,
  input         io_input_valid_1021,
  input         io_input_valid_1022,
  input         io_input_valid_1023,
  input         io_iormac_0,
  input         io_iormac_1,
  input         io_iormac_2,
  input         io_iormac_3,
  input         io_iormac_4,
  input         io_iormac_5,
  input         io_iormac_6,
  input         io_iormac_7,
  input         io_iormac_8,
  input         io_iormac_9,
  input         io_iormac_10,
  input         io_iormac_11,
  input         io_iormac_12,
  input         io_iormac_13,
  input         io_iormac_14,
  input         io_iormac_15,
  input         io_iormac_16,
  input         io_iormac_17,
  input         io_iormac_18,
  input         io_iormac_19,
  input         io_iormac_20,
  input         io_iormac_21,
  input         io_iormac_22,
  input         io_iormac_23,
  input         io_iormac_24,
  input         io_iormac_25,
  input         io_iormac_26,
  input         io_iormac_27,
  input         io_iormac_28,
  input         io_iormac_29,
  input         io_iormac_30,
  input         io_iormac_31,
  input         io_iormac_32,
  input         io_iormac_33,
  input         io_iormac_34,
  input         io_iormac_35,
  input         io_iormac_36,
  input         io_iormac_37,
  input         io_iormac_38,
  input         io_iormac_39,
  input         io_iormac_40,
  input         io_iormac_41,
  input         io_iormac_42,
  input         io_iormac_43,
  input         io_iormac_44,
  input         io_iormac_45,
  input         io_iormac_46,
  input         io_iormac_47,
  input         io_iormac_48,
  input         io_iormac_49,
  input         io_iormac_50,
  input         io_iormac_51,
  input         io_iormac_52,
  input         io_iormac_53,
  input         io_iormac_54,
  input         io_iormac_55,
  input         io_iormac_56,
  input         io_iormac_57,
  input         io_iormac_58,
  input         io_iormac_59,
  input         io_iormac_60,
  input         io_iormac_61,
  input         io_iormac_62,
  input         io_iormac_63,
  input         io_iormac_64,
  input         io_iormac_65,
  input         io_iormac_66,
  input         io_iormac_67,
  input         io_iormac_68,
  input         io_iormac_69,
  input         io_iormac_70,
  input         io_iormac_71,
  input         io_iormac_72,
  input         io_iormac_73,
  input         io_iormac_74,
  input         io_iormac_75,
  input         io_iormac_76,
  input         io_iormac_77,
  input         io_iormac_78,
  input         io_iormac_79,
  input         io_iormac_80,
  input         io_iormac_81,
  input         io_iormac_82,
  input         io_iormac_83,
  input         io_iormac_84,
  input         io_iormac_85,
  input         io_iormac_86,
  input         io_iormac_87,
  input         io_iormac_88,
  input         io_iormac_89,
  input         io_iormac_90,
  input         io_iormac_91,
  input         io_iormac_92,
  input         io_iormac_93,
  input         io_iormac_94,
  input         io_iormac_95,
  input         io_iormac_96,
  input         io_iormac_97,
  input         io_iormac_98,
  input         io_iormac_99,
  input         io_iormac_100,
  input         io_iormac_101,
  input         io_iormac_102,
  input         io_iormac_103,
  input         io_iormac_104,
  input         io_iormac_105,
  input         io_iormac_106,
  input         io_iormac_107,
  input         io_iormac_108,
  input         io_iormac_109,
  input         io_iormac_110,
  input         io_iormac_111,
  input         io_iormac_112,
  input         io_iormac_113,
  input         io_iormac_114,
  input         io_iormac_115,
  input         io_iormac_116,
  input         io_iormac_117,
  input         io_iormac_118,
  input         io_iormac_119,
  input         io_iormac_120,
  input         io_iormac_121,
  input         io_iormac_122,
  input         io_iormac_123,
  input         io_iormac_124,
  input         io_iormac_125,
  input         io_iormac_126,
  input         io_iormac_127,
  input         io_iormac_128,
  input         io_iormac_129,
  input         io_iormac_130,
  input         io_iormac_131,
  input         io_iormac_132,
  input         io_iormac_133,
  input         io_iormac_134,
  input         io_iormac_135,
  input         io_iormac_136,
  input         io_iormac_137,
  input         io_iormac_138,
  input         io_iormac_139,
  input         io_iormac_140,
  input         io_iormac_141,
  input         io_iormac_142,
  input         io_iormac_143,
  input         io_iormac_144,
  input         io_iormac_145,
  input         io_iormac_146,
  input         io_iormac_147,
  input         io_iormac_148,
  input         io_iormac_149,
  input         io_iormac_150,
  input         io_iormac_151,
  input         io_iormac_152,
  input         io_iormac_153,
  input         io_iormac_154,
  input         io_iormac_155,
  input         io_iormac_156,
  input         io_iormac_157,
  input         io_iormac_158,
  input         io_iormac_159,
  input         io_iormac_160,
  input         io_iormac_161,
  input         io_iormac_162,
  input         io_iormac_163,
  input         io_iormac_164,
  input         io_iormac_165,
  input         io_iormac_166,
  input         io_iormac_167,
  input         io_iormac_168,
  input         io_iormac_169,
  input         io_iormac_170,
  input         io_iormac_171,
  input         io_iormac_172,
  input         io_iormac_173,
  input         io_iormac_174,
  input         io_iormac_175,
  input         io_iormac_176,
  input         io_iormac_177,
  input         io_iormac_178,
  input         io_iormac_179,
  input         io_iormac_180,
  input         io_iormac_181,
  input         io_iormac_182,
  input         io_iormac_183,
  input         io_iormac_184,
  input         io_iormac_185,
  input         io_iormac_186,
  input         io_iormac_187,
  input         io_iormac_188,
  input         io_iormac_189,
  input         io_iormac_190,
  input         io_iormac_191,
  input         io_iormac_192,
  input         io_iormac_193,
  input         io_iormac_194,
  input         io_iormac_195,
  input         io_iormac_196,
  input         io_iormac_197,
  input         io_iormac_198,
  input         io_iormac_199,
  input         io_iormac_200,
  input         io_iormac_201,
  input         io_iormac_202,
  input         io_iormac_203,
  input         io_iormac_204,
  input         io_iormac_205,
  input         io_iormac_206,
  input         io_iormac_207,
  input         io_iormac_208,
  input         io_iormac_209,
  input         io_iormac_210,
  input         io_iormac_211,
  input         io_iormac_212,
  input         io_iormac_213,
  input         io_iormac_214,
  input         io_iormac_215,
  input         io_iormac_216,
  input         io_iormac_217,
  input         io_iormac_218,
  input         io_iormac_219,
  input         io_iormac_220,
  input         io_iormac_221,
  input         io_iormac_222,
  input         io_iormac_223,
  input         io_iormac_224,
  input         io_iormac_225,
  input         io_iormac_226,
  input         io_iormac_227,
  input         io_iormac_228,
  input         io_iormac_229,
  input         io_iormac_230,
  input         io_iormac_231,
  input         io_iormac_232,
  input         io_iormac_233,
  input         io_iormac_234,
  input         io_iormac_235,
  input         io_iormac_236,
  input         io_iormac_237,
  input         io_iormac_238,
  input         io_iormac_239,
  input         io_iormac_240,
  input         io_iormac_241,
  input         io_iormac_242,
  input         io_iormac_243,
  input         io_iormac_244,
  input         io_iormac_245,
  input         io_iormac_246,
  input         io_iormac_247,
  input         io_iormac_248,
  input         io_iormac_249,
  input         io_iormac_250,
  input         io_iormac_251,
  input         io_iormac_252,
  input         io_iormac_253,
  input         io_iormac_254,
  input         io_iormac_255,
  input         io_iormac_256,
  input         io_iormac_257,
  input         io_iormac_258,
  input         io_iormac_259,
  input         io_iormac_260,
  input         io_iormac_261,
  input         io_iormac_262,
  input         io_iormac_263,
  input         io_iormac_264,
  input         io_iormac_265,
  input         io_iormac_266,
  input         io_iormac_267,
  input         io_iormac_268,
  input         io_iormac_269,
  input         io_iormac_270,
  input         io_iormac_271,
  input         io_iormac_272,
  input         io_iormac_273,
  input         io_iormac_274,
  input         io_iormac_275,
  input         io_iormac_276,
  input         io_iormac_277,
  input         io_iormac_278,
  input         io_iormac_279,
  input         io_iormac_280,
  input         io_iormac_281,
  input         io_iormac_282,
  input         io_iormac_283,
  input         io_iormac_284,
  input         io_iormac_285,
  input         io_iormac_286,
  input         io_iormac_287,
  input         io_iormac_288,
  input         io_iormac_289,
  input         io_iormac_290,
  input         io_iormac_291,
  input         io_iormac_292,
  input         io_iormac_293,
  input         io_iormac_294,
  input         io_iormac_295,
  input         io_iormac_296,
  input         io_iormac_297,
  input         io_iormac_298,
  input         io_iormac_299,
  input         io_iormac_300,
  input         io_iormac_301,
  input         io_iormac_302,
  input         io_iormac_303,
  input         io_iormac_304,
  input         io_iormac_305,
  input         io_iormac_306,
  input         io_iormac_307,
  input         io_iormac_308,
  input         io_iormac_309,
  input         io_iormac_310,
  input         io_iormac_311,
  input         io_iormac_312,
  input         io_iormac_313,
  input         io_iormac_314,
  input         io_iormac_315,
  input         io_iormac_316,
  input         io_iormac_317,
  input         io_iormac_318,
  input         io_iormac_319,
  input         io_iormac_320,
  input         io_iormac_321,
  input         io_iormac_322,
  input         io_iormac_323,
  input         io_iormac_324,
  input         io_iormac_325,
  input         io_iormac_326,
  input         io_iormac_327,
  input         io_iormac_328,
  input         io_iormac_329,
  input         io_iormac_330,
  input         io_iormac_331,
  input         io_iormac_332,
  input         io_iormac_333,
  input         io_iormac_334,
  input         io_iormac_335,
  input         io_iormac_336,
  input         io_iormac_337,
  input         io_iormac_338,
  input         io_iormac_339,
  input         io_iormac_340,
  input         io_iormac_341,
  input         io_iormac_342,
  input         io_iormac_343,
  input         io_iormac_344,
  input         io_iormac_345,
  input         io_iormac_346,
  input         io_iormac_347,
  input         io_iormac_348,
  input         io_iormac_349,
  input         io_iormac_350,
  input         io_iormac_351,
  input         io_iormac_352,
  input         io_iormac_353,
  input         io_iormac_354,
  input         io_iormac_355,
  input         io_iormac_356,
  input         io_iormac_357,
  input         io_iormac_358,
  input         io_iormac_359,
  input         io_iormac_360,
  input         io_iormac_361,
  input         io_iormac_362,
  input         io_iormac_363,
  input         io_iormac_364,
  input         io_iormac_365,
  input         io_iormac_366,
  input         io_iormac_367,
  input         io_iormac_368,
  input         io_iormac_369,
  input         io_iormac_370,
  input         io_iormac_371,
  input         io_iormac_372,
  input         io_iormac_373,
  input         io_iormac_374,
  input         io_iormac_375,
  input         io_iormac_376,
  input         io_iormac_377,
  input         io_iormac_378,
  input         io_iormac_379,
  input         io_iormac_380,
  input         io_iormac_381,
  input         io_iormac_382,
  input         io_iormac_383,
  input         io_iormac_384,
  input         io_iormac_385,
  input         io_iormac_386,
  input         io_iormac_387,
  input         io_iormac_388,
  input         io_iormac_389,
  input         io_iormac_390,
  input         io_iormac_391,
  input         io_iormac_392,
  input         io_iormac_393,
  input         io_iormac_394,
  input         io_iormac_395,
  input         io_iormac_396,
  input         io_iormac_397,
  input         io_iormac_398,
  input         io_iormac_399,
  input         io_iormac_400,
  input         io_iormac_401,
  input         io_iormac_402,
  input         io_iormac_403,
  input         io_iormac_404,
  input         io_iormac_405,
  input         io_iormac_406,
  input         io_iormac_407,
  input         io_iormac_408,
  input         io_iormac_409,
  input         io_iormac_410,
  input         io_iormac_411,
  input         io_iormac_412,
  input         io_iormac_413,
  input         io_iormac_414,
  input         io_iormac_415,
  input         io_iormac_416,
  input         io_iormac_417,
  input         io_iormac_418,
  input         io_iormac_419,
  input         io_iormac_420,
  input         io_iormac_421,
  input         io_iormac_422,
  input         io_iormac_423,
  input         io_iormac_424,
  input         io_iormac_425,
  input         io_iormac_426,
  input         io_iormac_427,
  input         io_iormac_428,
  input         io_iormac_429,
  input         io_iormac_430,
  input         io_iormac_431,
  input         io_iormac_432,
  input         io_iormac_433,
  input         io_iormac_434,
  input         io_iormac_435,
  input         io_iormac_436,
  input         io_iormac_437,
  input         io_iormac_438,
  input         io_iormac_439,
  input         io_iormac_440,
  input         io_iormac_441,
  input         io_iormac_442,
  input         io_iormac_443,
  input         io_iormac_444,
  input         io_iormac_445,
  input         io_iormac_446,
  input         io_iormac_447,
  input         io_iormac_448,
  input         io_iormac_449,
  input         io_iormac_450,
  input         io_iormac_451,
  input         io_iormac_452,
  input         io_iormac_453,
  input         io_iormac_454,
  input         io_iormac_455,
  input         io_iormac_456,
  input         io_iormac_457,
  input         io_iormac_458,
  input         io_iormac_459,
  input         io_iormac_460,
  input         io_iormac_461,
  input         io_iormac_462,
  input         io_iormac_463,
  input         io_iormac_464,
  input         io_iormac_465,
  input         io_iormac_466,
  input         io_iormac_467,
  input         io_iormac_468,
  input         io_iormac_469,
  input         io_iormac_470,
  input         io_iormac_471,
  input         io_iormac_472,
  input         io_iormac_473,
  input         io_iormac_474,
  input         io_iormac_475,
  input         io_iormac_476,
  input         io_iormac_477,
  input         io_iormac_478,
  input         io_iormac_479,
  input         io_iormac_480,
  input         io_iormac_481,
  input         io_iormac_482,
  input         io_iormac_483,
  input         io_iormac_484,
  input         io_iormac_485,
  input         io_iormac_486,
  input         io_iormac_487,
  input         io_iormac_488,
  input         io_iormac_489,
  input         io_iormac_490,
  input         io_iormac_491,
  input         io_iormac_492,
  input         io_iormac_493,
  input         io_iormac_494,
  input         io_iormac_495,
  input         io_iormac_496,
  input         io_iormac_497,
  input         io_iormac_498,
  input         io_iormac_499,
  input         io_iormac_500,
  input         io_iormac_501,
  input         io_iormac_502,
  input         io_iormac_503,
  input         io_iormac_504,
  input         io_iormac_505,
  input         io_iormac_506,
  input         io_iormac_507,
  input         io_iormac_508,
  input         io_iormac_509,
  input         io_iormac_510,
  input         io_iormac_511,
  input         io_iormac_512,
  input         io_iormac_513,
  input         io_iormac_514,
  input         io_iormac_515,
  input         io_iormac_516,
  input         io_iormac_517,
  input         io_iormac_518,
  input         io_iormac_519,
  input         io_iormac_520,
  input         io_iormac_521,
  input         io_iormac_522,
  input         io_iormac_523,
  input         io_iormac_524,
  input         io_iormac_525,
  input         io_iormac_526,
  input         io_iormac_527,
  input         io_iormac_528,
  input         io_iormac_529,
  input         io_iormac_530,
  input         io_iormac_531,
  input         io_iormac_532,
  input         io_iormac_533,
  input         io_iormac_534,
  input         io_iormac_535,
  input         io_iormac_536,
  input         io_iormac_537,
  input         io_iormac_538,
  input         io_iormac_539,
  input         io_iormac_540,
  input         io_iormac_541,
  input         io_iormac_542,
  input         io_iormac_543,
  input         io_iormac_544,
  input         io_iormac_545,
  input         io_iormac_546,
  input         io_iormac_547,
  input         io_iormac_548,
  input         io_iormac_549,
  input         io_iormac_550,
  input         io_iormac_551,
  input         io_iormac_552,
  input         io_iormac_553,
  input         io_iormac_554,
  input         io_iormac_555,
  input         io_iormac_556,
  input         io_iormac_557,
  input         io_iormac_558,
  input         io_iormac_559,
  input         io_iormac_560,
  input         io_iormac_561,
  input         io_iormac_562,
  input         io_iormac_563,
  input         io_iormac_564,
  input         io_iormac_565,
  input         io_iormac_566,
  input         io_iormac_567,
  input         io_iormac_568,
  input         io_iormac_569,
  input         io_iormac_570,
  input         io_iormac_571,
  input         io_iormac_572,
  input         io_iormac_573,
  input         io_iormac_574,
  input         io_iormac_575,
  input         io_iormac_576,
  input         io_iormac_577,
  input         io_iormac_578,
  input         io_iormac_579,
  input         io_iormac_580,
  input         io_iormac_581,
  input         io_iormac_582,
  input         io_iormac_583,
  input         io_iormac_584,
  input         io_iormac_585,
  input         io_iormac_586,
  input         io_iormac_587,
  input         io_iormac_588,
  input         io_iormac_589,
  input         io_iormac_590,
  input         io_iormac_591,
  input         io_iormac_592,
  input         io_iormac_593,
  input         io_iormac_594,
  input         io_iormac_595,
  input         io_iormac_596,
  input         io_iormac_597,
  input         io_iormac_598,
  input         io_iormac_599,
  input         io_iormac_600,
  input         io_iormac_601,
  input         io_iormac_602,
  input         io_iormac_603,
  input         io_iormac_604,
  input         io_iormac_605,
  input         io_iormac_606,
  input         io_iormac_607,
  input         io_iormac_608,
  input         io_iormac_609,
  input         io_iormac_610,
  input         io_iormac_611,
  input         io_iormac_612,
  input         io_iormac_613,
  input         io_iormac_614,
  input         io_iormac_615,
  input         io_iormac_616,
  input         io_iormac_617,
  input         io_iormac_618,
  input         io_iormac_619,
  input         io_iormac_620,
  input         io_iormac_621,
  input         io_iormac_622,
  input         io_iormac_623,
  input         io_iormac_624,
  input         io_iormac_625,
  input         io_iormac_626,
  input         io_iormac_627,
  input         io_iormac_628,
  input         io_iormac_629,
  input         io_iormac_630,
  input         io_iormac_631,
  input         io_iormac_632,
  input         io_iormac_633,
  input         io_iormac_634,
  input         io_iormac_635,
  input         io_iormac_636,
  input         io_iormac_637,
  input         io_iormac_638,
  input         io_iormac_639,
  input         io_iormac_640,
  input         io_iormac_641,
  input         io_iormac_642,
  input         io_iormac_643,
  input         io_iormac_644,
  input         io_iormac_645,
  input         io_iormac_646,
  input         io_iormac_647,
  input         io_iormac_648,
  input         io_iormac_649,
  input         io_iormac_650,
  input         io_iormac_651,
  input         io_iormac_652,
  input         io_iormac_653,
  input         io_iormac_654,
  input         io_iormac_655,
  input         io_iormac_656,
  input         io_iormac_657,
  input         io_iormac_658,
  input         io_iormac_659,
  input         io_iormac_660,
  input         io_iormac_661,
  input         io_iormac_662,
  input         io_iormac_663,
  input         io_iormac_664,
  input         io_iormac_665,
  input         io_iormac_666,
  input         io_iormac_667,
  input         io_iormac_668,
  input         io_iormac_669,
  input         io_iormac_670,
  input         io_iormac_671,
  input         io_iormac_672,
  input         io_iormac_673,
  input         io_iormac_674,
  input         io_iormac_675,
  input         io_iormac_676,
  input         io_iormac_677,
  input         io_iormac_678,
  input         io_iormac_679,
  input         io_iormac_680,
  input         io_iormac_681,
  input         io_iormac_682,
  input         io_iormac_683,
  input         io_iormac_684,
  input         io_iormac_685,
  input         io_iormac_686,
  input         io_iormac_687,
  input         io_iormac_688,
  input         io_iormac_689,
  input         io_iormac_690,
  input         io_iormac_691,
  input         io_iormac_692,
  input         io_iormac_693,
  input         io_iormac_694,
  input         io_iormac_695,
  input         io_iormac_696,
  input         io_iormac_697,
  input         io_iormac_698,
  input         io_iormac_699,
  input         io_iormac_700,
  input         io_iormac_701,
  input         io_iormac_702,
  input         io_iormac_703,
  input         io_iormac_704,
  input         io_iormac_705,
  input         io_iormac_706,
  input         io_iormac_707,
  input         io_iormac_708,
  input         io_iormac_709,
  input         io_iormac_710,
  input         io_iormac_711,
  input         io_iormac_712,
  input         io_iormac_713,
  input         io_iormac_714,
  input         io_iormac_715,
  input         io_iormac_716,
  input         io_iormac_717,
  input         io_iormac_718,
  input         io_iormac_719,
  input         io_iormac_720,
  input         io_iormac_721,
  input         io_iormac_722,
  input         io_iormac_723,
  input         io_iormac_724,
  input         io_iormac_725,
  input         io_iormac_726,
  input         io_iormac_727,
  input         io_iormac_728,
  input         io_iormac_729,
  input         io_iormac_730,
  input         io_iormac_731,
  input         io_iormac_732,
  input         io_iormac_733,
  input         io_iormac_734,
  input         io_iormac_735,
  input         io_iormac_736,
  input         io_iormac_737,
  input         io_iormac_738,
  input         io_iormac_739,
  input         io_iormac_740,
  input         io_iormac_741,
  input         io_iormac_742,
  input         io_iormac_743,
  input         io_iormac_744,
  input         io_iormac_745,
  input         io_iormac_746,
  input         io_iormac_747,
  input         io_iormac_748,
  input         io_iormac_749,
  input         io_iormac_750,
  input         io_iormac_751,
  input         io_iormac_752,
  input         io_iormac_753,
  input         io_iormac_754,
  input         io_iormac_755,
  input         io_iormac_756,
  input         io_iormac_757,
  input         io_iormac_758,
  input         io_iormac_759,
  input         io_iormac_760,
  input         io_iormac_761,
  input         io_iormac_762,
  input         io_iormac_763,
  input         io_iormac_764,
  input         io_iormac_765,
  input         io_iormac_766,
  input         io_iormac_767,
  input         io_iormac_768,
  input         io_iormac_769,
  input         io_iormac_770,
  input         io_iormac_771,
  input         io_iormac_772,
  input         io_iormac_773,
  input         io_iormac_774,
  input         io_iormac_775,
  input         io_iormac_776,
  input         io_iormac_777,
  input         io_iormac_778,
  input         io_iormac_779,
  input         io_iormac_780,
  input         io_iormac_781,
  input         io_iormac_782,
  input         io_iormac_783,
  input         io_iormac_784,
  input         io_iormac_785,
  input         io_iormac_786,
  input         io_iormac_787,
  input         io_iormac_788,
  input         io_iormac_789,
  input         io_iormac_790,
  input         io_iormac_791,
  input         io_iormac_792,
  input         io_iormac_793,
  input         io_iormac_794,
  input         io_iormac_795,
  input         io_iormac_796,
  input         io_iormac_797,
  input         io_iormac_798,
  input         io_iormac_799,
  input         io_iormac_800,
  input         io_iormac_801,
  input         io_iormac_802,
  input         io_iormac_803,
  input         io_iormac_804,
  input         io_iormac_805,
  input         io_iormac_806,
  input         io_iormac_807,
  input         io_iormac_808,
  input         io_iormac_809,
  input         io_iormac_810,
  input         io_iormac_811,
  input         io_iormac_812,
  input         io_iormac_813,
  input         io_iormac_814,
  input         io_iormac_815,
  input         io_iormac_816,
  input         io_iormac_817,
  input         io_iormac_818,
  input         io_iormac_819,
  input         io_iormac_820,
  input         io_iormac_821,
  input         io_iormac_822,
  input         io_iormac_823,
  input         io_iormac_824,
  input         io_iormac_825,
  input         io_iormac_826,
  input         io_iormac_827,
  input         io_iormac_828,
  input         io_iormac_829,
  input         io_iormac_830,
  input         io_iormac_831,
  input         io_iormac_832,
  input         io_iormac_833,
  input         io_iormac_834,
  input         io_iormac_835,
  input         io_iormac_836,
  input         io_iormac_837,
  input         io_iormac_838,
  input         io_iormac_839,
  input         io_iormac_840,
  input         io_iormac_841,
  input         io_iormac_842,
  input         io_iormac_843,
  input         io_iormac_844,
  input         io_iormac_845,
  input         io_iormac_846,
  input         io_iormac_847,
  input         io_iormac_848,
  input         io_iormac_849,
  input         io_iormac_850,
  input         io_iormac_851,
  input         io_iormac_852,
  input         io_iormac_853,
  input         io_iormac_854,
  input         io_iormac_855,
  input         io_iormac_856,
  input         io_iormac_857,
  input         io_iormac_858,
  input         io_iormac_859,
  input         io_iormac_860,
  input         io_iormac_861,
  input         io_iormac_862,
  input         io_iormac_863,
  input         io_iormac_864,
  input         io_iormac_865,
  input         io_iormac_866,
  input         io_iormac_867,
  input         io_iormac_868,
  input         io_iormac_869,
  input         io_iormac_870,
  input         io_iormac_871,
  input         io_iormac_872,
  input         io_iormac_873,
  input         io_iormac_874,
  input         io_iormac_875,
  input         io_iormac_876,
  input         io_iormac_877,
  input         io_iormac_878,
  input         io_iormac_879,
  input         io_iormac_880,
  input         io_iormac_881,
  input         io_iormac_882,
  input         io_iormac_883,
  input         io_iormac_884,
  input         io_iormac_885,
  input         io_iormac_886,
  input         io_iormac_887,
  input         io_iormac_888,
  input         io_iormac_889,
  input         io_iormac_890,
  input         io_iormac_891,
  input         io_iormac_892,
  input         io_iormac_893,
  input         io_iormac_894,
  input         io_iormac_895,
  input         io_iormac_896,
  input         io_iormac_897,
  input         io_iormac_898,
  input         io_iormac_899,
  input         io_iormac_900,
  input         io_iormac_901,
  input         io_iormac_902,
  input         io_iormac_903,
  input         io_iormac_904,
  input         io_iormac_905,
  input         io_iormac_906,
  input         io_iormac_907,
  input         io_iormac_908,
  input         io_iormac_909,
  input         io_iormac_910,
  input         io_iormac_911,
  input         io_iormac_912,
  input         io_iormac_913,
  input         io_iormac_914,
  input         io_iormac_915,
  input         io_iormac_916,
  input         io_iormac_917,
  input         io_iormac_918,
  input         io_iormac_919,
  input         io_iormac_920,
  input         io_iormac_921,
  input         io_iormac_922,
  input         io_iormac_923,
  input         io_iormac_924,
  input         io_iormac_925,
  input         io_iormac_926,
  input         io_iormac_927,
  input         io_iormac_928,
  input         io_iormac_929,
  input         io_iormac_930,
  input         io_iormac_931,
  input         io_iormac_932,
  input         io_iormac_933,
  input         io_iormac_934,
  input         io_iormac_935,
  input         io_iormac_936,
  input         io_iormac_937,
  input         io_iormac_938,
  input         io_iormac_939,
  input         io_iormac_940,
  input         io_iormac_941,
  input         io_iormac_942,
  input         io_iormac_943,
  input         io_iormac_944,
  input         io_iormac_945,
  input         io_iormac_946,
  input         io_iormac_947,
  input         io_iormac_948,
  input         io_iormac_949,
  input         io_iormac_950,
  input         io_iormac_951,
  input         io_iormac_952,
  input         io_iormac_953,
  input         io_iormac_954,
  input         io_iormac_955,
  input         io_iormac_956,
  input         io_iormac_957,
  input         io_iormac_958,
  input         io_iormac_959,
  input         io_iormac_960,
  input         io_iormac_961,
  input         io_iormac_962,
  input         io_iormac_963,
  input         io_iormac_964,
  input         io_iormac_965,
  input         io_iormac_966,
  input         io_iormac_967,
  input         io_iormac_968,
  input         io_iormac_969,
  input         io_iormac_970,
  input         io_iormac_971,
  input         io_iormac_972,
  input         io_iormac_973,
  input         io_iormac_974,
  input         io_iormac_975,
  input         io_iormac_976,
  input         io_iormac_977,
  input         io_iormac_978,
  input         io_iormac_979,
  input         io_iormac_980,
  input         io_iormac_981,
  input         io_iormac_982,
  input         io_iormac_983,
  input         io_iormac_984,
  input         io_iormac_985,
  input         io_iormac_986,
  input         io_iormac_987,
  input         io_iormac_988,
  input         io_iormac_989,
  input         io_iormac_990,
  input         io_iormac_991,
  input         io_iormac_992,
  input         io_iormac_993,
  input         io_iormac_994,
  input         io_iormac_995,
  input         io_iormac_996,
  input         io_iormac_997,
  input         io_iormac_998,
  input         io_iormac_999,
  input         io_iormac_1000,
  input         io_iormac_1001,
  input         io_iormac_1002,
  input         io_iormac_1003,
  input         io_iormac_1004,
  input         io_iormac_1005,
  input         io_iormac_1006,
  input         io_iormac_1007,
  input         io_iormac_1008,
  input         io_iormac_1009,
  input         io_iormac_1010,
  input         io_iormac_1011,
  input         io_iormac_1012,
  input         io_iormac_1013,
  input         io_iormac_1014,
  input         io_iormac_1015,
  input         io_iormac_1016,
  input         io_iormac_1017,
  input         io_iormac_1018,
  input         io_iormac_1019,
  input         io_iormac_1020,
  input         io_iormac_1021,
  input         io_iormac_1022,
  input         io_iormac_1023,
  output [31:0] io_out_0,
  output [31:0] io_out_1,
  output [31:0] io_out_2,
  output [31:0] io_out_3,
  output [31:0] io_out_4,
  output [31:0] io_out_5,
  output [31:0] io_out_6,
  output [31:0] io_out_7,
  output [31:0] io_out_8,
  output [31:0] io_out_9,
  output [31:0] io_out_10,
  output [31:0] io_out_11,
  output [31:0] io_out_12,
  output [31:0] io_out_13,
  output [31:0] io_out_14,
  output [31:0] io_out_15,
  output [31:0] io_out_16,
  output [31:0] io_out_17,
  output [31:0] io_out_18,
  output [31:0] io_out_19,
  output [31:0] io_out_20,
  output [31:0] io_out_21,
  output [31:0] io_out_22,
  output [31:0] io_out_23,
  output [31:0] io_out_24,
  output [31:0] io_out_25,
  output [31:0] io_out_26,
  output [31:0] io_out_27,
  output [31:0] io_out_28,
  output [31:0] io_out_29,
  output [31:0] io_out_30,
  output [31:0] io_out_31,
  output [31:0] io_out_32,
  output [31:0] io_out_33,
  output [31:0] io_out_34,
  output [31:0] io_out_35,
  output [31:0] io_out_36,
  output [31:0] io_out_37,
  output [31:0] io_out_38,
  output [31:0] io_out_39,
  output [31:0] io_out_40,
  output [31:0] io_out_41,
  output [31:0] io_out_42,
  output [31:0] io_out_43,
  output [31:0] io_out_44,
  output [31:0] io_out_45,
  output [31:0] io_out_46,
  output [31:0] io_out_47,
  output [31:0] io_out_48,
  output [31:0] io_out_49,
  output [31:0] io_out_50,
  output [31:0] io_out_51,
  output [31:0] io_out_52,
  output [31:0] io_out_53,
  output [31:0] io_out_54,
  output [31:0] io_out_55,
  output [31:0] io_out_56,
  output [31:0] io_out_57,
  output [31:0] io_out_58,
  output [31:0] io_out_59,
  output [31:0] io_out_60,
  output [31:0] io_out_61,
  output [31:0] io_out_62,
  output [31:0] io_out_63,
  output [31:0] io_out_64,
  output [31:0] io_out_65,
  output [31:0] io_out_66,
  output [31:0] io_out_67,
  output [31:0] io_out_68,
  output [31:0] io_out_69,
  output [31:0] io_out_70,
  output [31:0] io_out_71,
  output [31:0] io_out_72,
  output [31:0] io_out_73,
  output [31:0] io_out_74,
  output [31:0] io_out_75,
  output [31:0] io_out_76,
  output [31:0] io_out_77,
  output [31:0] io_out_78,
  output [31:0] io_out_79,
  output [31:0] io_out_80,
  output [31:0] io_out_81,
  output [31:0] io_out_82,
  output [31:0] io_out_83,
  output [31:0] io_out_84,
  output [31:0] io_out_85,
  output [31:0] io_out_86,
  output [31:0] io_out_87,
  output [31:0] io_out_88,
  output [31:0] io_out_89,
  output [31:0] io_out_90,
  output [31:0] io_out_91,
  output [31:0] io_out_92,
  output [31:0] io_out_93,
  output [31:0] io_out_94,
  output [31:0] io_out_95,
  output [31:0] io_out_96,
  output [31:0] io_out_97,
  output [31:0] io_out_98,
  output [31:0] io_out_99,
  output [31:0] io_out_100,
  output [31:0] io_out_101,
  output [31:0] io_out_102,
  output [31:0] io_out_103,
  output [31:0] io_out_104,
  output [31:0] io_out_105,
  output [31:0] io_out_106,
  output [31:0] io_out_107,
  output [31:0] io_out_108,
  output [31:0] io_out_109,
  output [31:0] io_out_110,
  output [31:0] io_out_111,
  output [31:0] io_out_112,
  output [31:0] io_out_113,
  output [31:0] io_out_114,
  output [31:0] io_out_115,
  output [31:0] io_out_116,
  output [31:0] io_out_117,
  output [31:0] io_out_118,
  output [31:0] io_out_119,
  output [31:0] io_out_120,
  output [31:0] io_out_121,
  output [31:0] io_out_122,
  output [31:0] io_out_123,
  output [31:0] io_out_124,
  output [31:0] io_out_125,
  output [31:0] io_out_126,
  output [31:0] io_out_127,
  output [31:0] io_out_128,
  output [31:0] io_out_129,
  output [31:0] io_out_130,
  output [31:0] io_out_131,
  output [31:0] io_out_132,
  output [31:0] io_out_133,
  output [31:0] io_out_134,
  output [31:0] io_out_135,
  output [31:0] io_out_136,
  output [31:0] io_out_137,
  output [31:0] io_out_138,
  output [31:0] io_out_139,
  output [31:0] io_out_140,
  output [31:0] io_out_141,
  output [31:0] io_out_142,
  output [31:0] io_out_143,
  output [31:0] io_out_144,
  output [31:0] io_out_145,
  output [31:0] io_out_146,
  output [31:0] io_out_147,
  output [31:0] io_out_148,
  output [31:0] io_out_149,
  output [31:0] io_out_150,
  output [31:0] io_out_151,
  output [31:0] io_out_152,
  output [31:0] io_out_153,
  output [31:0] io_out_154,
  output [31:0] io_out_155,
  output [31:0] io_out_156,
  output [31:0] io_out_157,
  output [31:0] io_out_158,
  output [31:0] io_out_159,
  output [31:0] io_out_160,
  output [31:0] io_out_161,
  output [31:0] io_out_162,
  output [31:0] io_out_163,
  output [31:0] io_out_164,
  output [31:0] io_out_165,
  output [31:0] io_out_166,
  output [31:0] io_out_167,
  output [31:0] io_out_168,
  output [31:0] io_out_169,
  output [31:0] io_out_170,
  output [31:0] io_out_171,
  output [31:0] io_out_172,
  output [31:0] io_out_173,
  output [31:0] io_out_174,
  output [31:0] io_out_175,
  output [31:0] io_out_176,
  output [31:0] io_out_177,
  output [31:0] io_out_178,
  output [31:0] io_out_179,
  output [31:0] io_out_180,
  output [31:0] io_out_181,
  output [31:0] io_out_182,
  output [31:0] io_out_183,
  output [31:0] io_out_184,
  output [31:0] io_out_185,
  output [31:0] io_out_186,
  output [31:0] io_out_187,
  output [31:0] io_out_188,
  output [31:0] io_out_189,
  output [31:0] io_out_190,
  output [31:0] io_out_191,
  output [31:0] io_out_192,
  output [31:0] io_out_193,
  output [31:0] io_out_194,
  output [31:0] io_out_195,
  output [31:0] io_out_196,
  output [31:0] io_out_197,
  output [31:0] io_out_198,
  output [31:0] io_out_199,
  output [31:0] io_out_200,
  output [31:0] io_out_201,
  output [31:0] io_out_202,
  output [31:0] io_out_203,
  output [31:0] io_out_204,
  output [31:0] io_out_205,
  output [31:0] io_out_206,
  output [31:0] io_out_207,
  output [31:0] io_out_208,
  output [31:0] io_out_209,
  output [31:0] io_out_210,
  output [31:0] io_out_211,
  output [31:0] io_out_212,
  output [31:0] io_out_213,
  output [31:0] io_out_214,
  output [31:0] io_out_215,
  output [31:0] io_out_216,
  output [31:0] io_out_217,
  output [31:0] io_out_218,
  output [31:0] io_out_219,
  output [31:0] io_out_220,
  output [31:0] io_out_221,
  output [31:0] io_out_222,
  output [31:0] io_out_223,
  output [31:0] io_out_224,
  output [31:0] io_out_225,
  output [31:0] io_out_226,
  output [31:0] io_out_227,
  output [31:0] io_out_228,
  output [31:0] io_out_229,
  output [31:0] io_out_230,
  output [31:0] io_out_231,
  output [31:0] io_out_232,
  output [31:0] io_out_233,
  output [31:0] io_out_234,
  output [31:0] io_out_235,
  output [31:0] io_out_236,
  output [31:0] io_out_237,
  output [31:0] io_out_238,
  output [31:0] io_out_239,
  output [31:0] io_out_240,
  output [31:0] io_out_241,
  output [31:0] io_out_242,
  output [31:0] io_out_243,
  output [31:0] io_out_244,
  output [31:0] io_out_245,
  output [31:0] io_out_246,
  output [31:0] io_out_247,
  output [31:0] io_out_248,
  output [31:0] io_out_249,
  output [31:0] io_out_250,
  output [31:0] io_out_251,
  output [31:0] io_out_252,
  output [31:0] io_out_253,
  output [31:0] io_out_254,
  output [31:0] io_out_255,
  output [31:0] io_out_256,
  output [31:0] io_out_257,
  output [31:0] io_out_258,
  output [31:0] io_out_259,
  output [31:0] io_out_260,
  output [31:0] io_out_261,
  output [31:0] io_out_262,
  output [31:0] io_out_263,
  output [31:0] io_out_264,
  output [31:0] io_out_265,
  output [31:0] io_out_266,
  output [31:0] io_out_267,
  output [31:0] io_out_268,
  output [31:0] io_out_269,
  output [31:0] io_out_270,
  output [31:0] io_out_271,
  output [31:0] io_out_272,
  output [31:0] io_out_273,
  output [31:0] io_out_274,
  output [31:0] io_out_275,
  output [31:0] io_out_276,
  output [31:0] io_out_277,
  output [31:0] io_out_278,
  output [31:0] io_out_279,
  output [31:0] io_out_280,
  output [31:0] io_out_281,
  output [31:0] io_out_282,
  output [31:0] io_out_283,
  output [31:0] io_out_284,
  output [31:0] io_out_285,
  output [31:0] io_out_286,
  output [31:0] io_out_287,
  output [31:0] io_out_288,
  output [31:0] io_out_289,
  output [31:0] io_out_290,
  output [31:0] io_out_291,
  output [31:0] io_out_292,
  output [31:0] io_out_293,
  output [31:0] io_out_294,
  output [31:0] io_out_295,
  output [31:0] io_out_296,
  output [31:0] io_out_297,
  output [31:0] io_out_298,
  output [31:0] io_out_299,
  output [31:0] io_out_300,
  output [31:0] io_out_301,
  output [31:0] io_out_302,
  output [31:0] io_out_303,
  output [31:0] io_out_304,
  output [31:0] io_out_305,
  output [31:0] io_out_306,
  output [31:0] io_out_307,
  output [31:0] io_out_308,
  output [31:0] io_out_309,
  output [31:0] io_out_310,
  output [31:0] io_out_311,
  output [31:0] io_out_312,
  output [31:0] io_out_313,
  output [31:0] io_out_314,
  output [31:0] io_out_315,
  output [31:0] io_out_316,
  output [31:0] io_out_317,
  output [31:0] io_out_318,
  output [31:0] io_out_319,
  output [31:0] io_out_320,
  output [31:0] io_out_321,
  output [31:0] io_out_322,
  output [31:0] io_out_323,
  output [31:0] io_out_324,
  output [31:0] io_out_325,
  output [31:0] io_out_326,
  output [31:0] io_out_327,
  output [31:0] io_out_328,
  output [31:0] io_out_329,
  output [31:0] io_out_330,
  output [31:0] io_out_331,
  output [31:0] io_out_332,
  output [31:0] io_out_333,
  output [31:0] io_out_334,
  output [31:0] io_out_335,
  output [31:0] io_out_336,
  output [31:0] io_out_337,
  output [31:0] io_out_338,
  output [31:0] io_out_339,
  output [31:0] io_out_340,
  output [31:0] io_out_341,
  output [31:0] io_out_342,
  output [31:0] io_out_343,
  output [31:0] io_out_344,
  output [31:0] io_out_345,
  output [31:0] io_out_346,
  output [31:0] io_out_347,
  output [31:0] io_out_348,
  output [31:0] io_out_349,
  output [31:0] io_out_350,
  output [31:0] io_out_351,
  output [31:0] io_out_352,
  output [31:0] io_out_353,
  output [31:0] io_out_354,
  output [31:0] io_out_355,
  output [31:0] io_out_356,
  output [31:0] io_out_357,
  output [31:0] io_out_358,
  output [31:0] io_out_359,
  output [31:0] io_out_360,
  output [31:0] io_out_361,
  output [31:0] io_out_362,
  output [31:0] io_out_363,
  output [31:0] io_out_364,
  output [31:0] io_out_365,
  output [31:0] io_out_366,
  output [31:0] io_out_367,
  output [31:0] io_out_368,
  output [31:0] io_out_369,
  output [31:0] io_out_370,
  output [31:0] io_out_371,
  output [31:0] io_out_372,
  output [31:0] io_out_373,
  output [31:0] io_out_374,
  output [31:0] io_out_375,
  output [31:0] io_out_376,
  output [31:0] io_out_377,
  output [31:0] io_out_378,
  output [31:0] io_out_379,
  output [31:0] io_out_380,
  output [31:0] io_out_381,
  output [31:0] io_out_382,
  output [31:0] io_out_383,
  output [31:0] io_out_384,
  output [31:0] io_out_385,
  output [31:0] io_out_386,
  output [31:0] io_out_387,
  output [31:0] io_out_388,
  output [31:0] io_out_389,
  output [31:0] io_out_390,
  output [31:0] io_out_391,
  output [31:0] io_out_392,
  output [31:0] io_out_393,
  output [31:0] io_out_394,
  output [31:0] io_out_395,
  output [31:0] io_out_396,
  output [31:0] io_out_397,
  output [31:0] io_out_398,
  output [31:0] io_out_399,
  output [31:0] io_out_400,
  output [31:0] io_out_401,
  output [31:0] io_out_402,
  output [31:0] io_out_403,
  output [31:0] io_out_404,
  output [31:0] io_out_405,
  output [31:0] io_out_406,
  output [31:0] io_out_407,
  output [31:0] io_out_408,
  output [31:0] io_out_409,
  output [31:0] io_out_410,
  output [31:0] io_out_411,
  output [31:0] io_out_412,
  output [31:0] io_out_413,
  output [31:0] io_out_414,
  output [31:0] io_out_415,
  output [31:0] io_out_416,
  output [31:0] io_out_417,
  output [31:0] io_out_418,
  output [31:0] io_out_419,
  output [31:0] io_out_420,
  output [31:0] io_out_421,
  output [31:0] io_out_422,
  output [31:0] io_out_423,
  output [31:0] io_out_424,
  output [31:0] io_out_425,
  output [31:0] io_out_426,
  output [31:0] io_out_427,
  output [31:0] io_out_428,
  output [31:0] io_out_429,
  output [31:0] io_out_430,
  output [31:0] io_out_431,
  output [31:0] io_out_432,
  output [31:0] io_out_433,
  output [31:0] io_out_434,
  output [31:0] io_out_435,
  output [31:0] io_out_436,
  output [31:0] io_out_437,
  output [31:0] io_out_438,
  output [31:0] io_out_439,
  output [31:0] io_out_440,
  output [31:0] io_out_441,
  output [31:0] io_out_442,
  output [31:0] io_out_443,
  output [31:0] io_out_444,
  output [31:0] io_out_445,
  output [31:0] io_out_446,
  output [31:0] io_out_447,
  output [31:0] io_out_448,
  output [31:0] io_out_449,
  output [31:0] io_out_450,
  output [31:0] io_out_451,
  output [31:0] io_out_452,
  output [31:0] io_out_453,
  output [31:0] io_out_454,
  output [31:0] io_out_455,
  output [31:0] io_out_456,
  output [31:0] io_out_457,
  output [31:0] io_out_458,
  output [31:0] io_out_459,
  output [31:0] io_out_460,
  output [31:0] io_out_461,
  output [31:0] io_out_462,
  output [31:0] io_out_463,
  output [31:0] io_out_464,
  output [31:0] io_out_465,
  output [31:0] io_out_466,
  output [31:0] io_out_467,
  output [31:0] io_out_468,
  output [31:0] io_out_469,
  output [31:0] io_out_470,
  output [31:0] io_out_471,
  output [31:0] io_out_472,
  output [31:0] io_out_473,
  output [31:0] io_out_474,
  output [31:0] io_out_475,
  output [31:0] io_out_476,
  output [31:0] io_out_477,
  output [31:0] io_out_478,
  output [31:0] io_out_479,
  output [31:0] io_out_480,
  output [31:0] io_out_481,
  output [31:0] io_out_482,
  output [31:0] io_out_483,
  output [31:0] io_out_484,
  output [31:0] io_out_485,
  output [31:0] io_out_486,
  output [31:0] io_out_487,
  output [31:0] io_out_488,
  output [31:0] io_out_489,
  output [31:0] io_out_490,
  output [31:0] io_out_491,
  output [31:0] io_out_492,
  output [31:0] io_out_493,
  output [31:0] io_out_494,
  output [31:0] io_out_495,
  output [31:0] io_out_496,
  output [31:0] io_out_497,
  output [31:0] io_out_498,
  output [31:0] io_out_499,
  output [31:0] io_out_500,
  output [31:0] io_out_501,
  output [31:0] io_out_502,
  output [31:0] io_out_503,
  output [31:0] io_out_504,
  output [31:0] io_out_505,
  output [31:0] io_out_506,
  output [31:0] io_out_507,
  output [31:0] io_out_508,
  output [31:0] io_out_509,
  output [31:0] io_out_510,
  output [31:0] io_out_511,
  output [31:0] io_out_512,
  output [31:0] io_out_513,
  output [31:0] io_out_514,
  output [31:0] io_out_515,
  output [31:0] io_out_516,
  output [31:0] io_out_517,
  output [31:0] io_out_518,
  output [31:0] io_out_519,
  output [31:0] io_out_520,
  output [31:0] io_out_521,
  output [31:0] io_out_522,
  output [31:0] io_out_523,
  output [31:0] io_out_524,
  output [31:0] io_out_525,
  output [31:0] io_out_526,
  output [31:0] io_out_527,
  output [31:0] io_out_528,
  output [31:0] io_out_529,
  output [31:0] io_out_530,
  output [31:0] io_out_531,
  output [31:0] io_out_532,
  output [31:0] io_out_533,
  output [31:0] io_out_534,
  output [31:0] io_out_535,
  output [31:0] io_out_536,
  output [31:0] io_out_537,
  output [31:0] io_out_538,
  output [31:0] io_out_539,
  output [31:0] io_out_540,
  output [31:0] io_out_541,
  output [31:0] io_out_542,
  output [31:0] io_out_543,
  output [31:0] io_out_544,
  output [31:0] io_out_545,
  output [31:0] io_out_546,
  output [31:0] io_out_547,
  output [31:0] io_out_548,
  output [31:0] io_out_549,
  output [31:0] io_out_550,
  output [31:0] io_out_551,
  output [31:0] io_out_552,
  output [31:0] io_out_553,
  output [31:0] io_out_554,
  output [31:0] io_out_555,
  output [31:0] io_out_556,
  output [31:0] io_out_557,
  output [31:0] io_out_558,
  output [31:0] io_out_559,
  output [31:0] io_out_560,
  output [31:0] io_out_561,
  output [31:0] io_out_562,
  output [31:0] io_out_563,
  output [31:0] io_out_564,
  output [31:0] io_out_565,
  output [31:0] io_out_566,
  output [31:0] io_out_567,
  output [31:0] io_out_568,
  output [31:0] io_out_569,
  output [31:0] io_out_570,
  output [31:0] io_out_571,
  output [31:0] io_out_572,
  output [31:0] io_out_573,
  output [31:0] io_out_574,
  output [31:0] io_out_575,
  output [31:0] io_out_576,
  output [31:0] io_out_577,
  output [31:0] io_out_578,
  output [31:0] io_out_579,
  output [31:0] io_out_580,
  output [31:0] io_out_581,
  output [31:0] io_out_582,
  output [31:0] io_out_583,
  output [31:0] io_out_584,
  output [31:0] io_out_585,
  output [31:0] io_out_586,
  output [31:0] io_out_587,
  output [31:0] io_out_588,
  output [31:0] io_out_589,
  output [31:0] io_out_590,
  output [31:0] io_out_591,
  output [31:0] io_out_592,
  output [31:0] io_out_593,
  output [31:0] io_out_594,
  output [31:0] io_out_595,
  output [31:0] io_out_596,
  output [31:0] io_out_597,
  output [31:0] io_out_598,
  output [31:0] io_out_599,
  output [31:0] io_out_600,
  output [31:0] io_out_601,
  output [31:0] io_out_602,
  output [31:0] io_out_603,
  output [31:0] io_out_604,
  output [31:0] io_out_605,
  output [31:0] io_out_606,
  output [31:0] io_out_607,
  output [31:0] io_out_608,
  output [31:0] io_out_609,
  output [31:0] io_out_610,
  output [31:0] io_out_611,
  output [31:0] io_out_612,
  output [31:0] io_out_613,
  output [31:0] io_out_614,
  output [31:0] io_out_615,
  output [31:0] io_out_616,
  output [31:0] io_out_617,
  output [31:0] io_out_618,
  output [31:0] io_out_619,
  output [31:0] io_out_620,
  output [31:0] io_out_621,
  output [31:0] io_out_622,
  output [31:0] io_out_623,
  output [31:0] io_out_624,
  output [31:0] io_out_625,
  output [31:0] io_out_626,
  output [31:0] io_out_627,
  output [31:0] io_out_628,
  output [31:0] io_out_629,
  output [31:0] io_out_630,
  output [31:0] io_out_631,
  output [31:0] io_out_632,
  output [31:0] io_out_633,
  output [31:0] io_out_634,
  output [31:0] io_out_635,
  output [31:0] io_out_636,
  output [31:0] io_out_637,
  output [31:0] io_out_638,
  output [31:0] io_out_639,
  output [31:0] io_out_640,
  output [31:0] io_out_641,
  output [31:0] io_out_642,
  output [31:0] io_out_643,
  output [31:0] io_out_644,
  output [31:0] io_out_645,
  output [31:0] io_out_646,
  output [31:0] io_out_647,
  output [31:0] io_out_648,
  output [31:0] io_out_649,
  output [31:0] io_out_650,
  output [31:0] io_out_651,
  output [31:0] io_out_652,
  output [31:0] io_out_653,
  output [31:0] io_out_654,
  output [31:0] io_out_655,
  output [31:0] io_out_656,
  output [31:0] io_out_657,
  output [31:0] io_out_658,
  output [31:0] io_out_659,
  output [31:0] io_out_660,
  output [31:0] io_out_661,
  output [31:0] io_out_662,
  output [31:0] io_out_663,
  output [31:0] io_out_664,
  output [31:0] io_out_665,
  output [31:0] io_out_666,
  output [31:0] io_out_667,
  output [31:0] io_out_668,
  output [31:0] io_out_669,
  output [31:0] io_out_670,
  output [31:0] io_out_671,
  output [31:0] io_out_672,
  output [31:0] io_out_673,
  output [31:0] io_out_674,
  output [31:0] io_out_675,
  output [31:0] io_out_676,
  output [31:0] io_out_677,
  output [31:0] io_out_678,
  output [31:0] io_out_679,
  output [31:0] io_out_680,
  output [31:0] io_out_681,
  output [31:0] io_out_682,
  output [31:0] io_out_683,
  output [31:0] io_out_684,
  output [31:0] io_out_685,
  output [31:0] io_out_686,
  output [31:0] io_out_687,
  output [31:0] io_out_688,
  output [31:0] io_out_689,
  output [31:0] io_out_690,
  output [31:0] io_out_691,
  output [31:0] io_out_692,
  output [31:0] io_out_693,
  output [31:0] io_out_694,
  output [31:0] io_out_695,
  output [31:0] io_out_696,
  output [31:0] io_out_697,
  output [31:0] io_out_698,
  output [31:0] io_out_699,
  output [31:0] io_out_700,
  output [31:0] io_out_701,
  output [31:0] io_out_702,
  output [31:0] io_out_703,
  output [31:0] io_out_704,
  output [31:0] io_out_705,
  output [31:0] io_out_706,
  output [31:0] io_out_707,
  output [31:0] io_out_708,
  output [31:0] io_out_709,
  output [31:0] io_out_710,
  output [31:0] io_out_711,
  output [31:0] io_out_712,
  output [31:0] io_out_713,
  output [31:0] io_out_714,
  output [31:0] io_out_715,
  output [31:0] io_out_716,
  output [31:0] io_out_717,
  output [31:0] io_out_718,
  output [31:0] io_out_719,
  output [31:0] io_out_720,
  output [31:0] io_out_721,
  output [31:0] io_out_722,
  output [31:0] io_out_723,
  output [31:0] io_out_724,
  output [31:0] io_out_725,
  output [31:0] io_out_726,
  output [31:0] io_out_727,
  output [31:0] io_out_728,
  output [31:0] io_out_729,
  output [31:0] io_out_730,
  output [31:0] io_out_731,
  output [31:0] io_out_732,
  output [31:0] io_out_733,
  output [31:0] io_out_734,
  output [31:0] io_out_735,
  output [31:0] io_out_736,
  output [31:0] io_out_737,
  output [31:0] io_out_738,
  output [31:0] io_out_739,
  output [31:0] io_out_740,
  output [31:0] io_out_741,
  output [31:0] io_out_742,
  output [31:0] io_out_743,
  output [31:0] io_out_744,
  output [31:0] io_out_745,
  output [31:0] io_out_746,
  output [31:0] io_out_747,
  output [31:0] io_out_748,
  output [31:0] io_out_749,
  output [31:0] io_out_750,
  output [31:0] io_out_751,
  output [31:0] io_out_752,
  output [31:0] io_out_753,
  output [31:0] io_out_754,
  output [31:0] io_out_755,
  output [31:0] io_out_756,
  output [31:0] io_out_757,
  output [31:0] io_out_758,
  output [31:0] io_out_759,
  output [31:0] io_out_760,
  output [31:0] io_out_761,
  output [31:0] io_out_762,
  output [31:0] io_out_763,
  output [31:0] io_out_764,
  output [31:0] io_out_765,
  output [31:0] io_out_766,
  output [31:0] io_out_767,
  output [31:0] io_out_768,
  output [31:0] io_out_769,
  output [31:0] io_out_770,
  output [31:0] io_out_771,
  output [31:0] io_out_772,
  output [31:0] io_out_773,
  output [31:0] io_out_774,
  output [31:0] io_out_775,
  output [31:0] io_out_776,
  output [31:0] io_out_777,
  output [31:0] io_out_778,
  output [31:0] io_out_779,
  output [31:0] io_out_780,
  output [31:0] io_out_781,
  output [31:0] io_out_782,
  output [31:0] io_out_783,
  output [31:0] io_out_784,
  output [31:0] io_out_785,
  output [31:0] io_out_786,
  output [31:0] io_out_787,
  output [31:0] io_out_788,
  output [31:0] io_out_789,
  output [31:0] io_out_790,
  output [31:0] io_out_791,
  output [31:0] io_out_792,
  output [31:0] io_out_793,
  output [31:0] io_out_794,
  output [31:0] io_out_795,
  output [31:0] io_out_796,
  output [31:0] io_out_797,
  output [31:0] io_out_798,
  output [31:0] io_out_799,
  output [31:0] io_out_800,
  output [31:0] io_out_801,
  output [31:0] io_out_802,
  output [31:0] io_out_803,
  output [31:0] io_out_804,
  output [31:0] io_out_805,
  output [31:0] io_out_806,
  output [31:0] io_out_807,
  output [31:0] io_out_808,
  output [31:0] io_out_809,
  output [31:0] io_out_810,
  output [31:0] io_out_811,
  output [31:0] io_out_812,
  output [31:0] io_out_813,
  output [31:0] io_out_814,
  output [31:0] io_out_815,
  output [31:0] io_out_816,
  output [31:0] io_out_817,
  output [31:0] io_out_818,
  output [31:0] io_out_819,
  output [31:0] io_out_820,
  output [31:0] io_out_821,
  output [31:0] io_out_822,
  output [31:0] io_out_823,
  output [31:0] io_out_824,
  output [31:0] io_out_825,
  output [31:0] io_out_826,
  output [31:0] io_out_827,
  output [31:0] io_out_828,
  output [31:0] io_out_829,
  output [31:0] io_out_830,
  output [31:0] io_out_831,
  output [31:0] io_out_832,
  output [31:0] io_out_833,
  output [31:0] io_out_834,
  output [31:0] io_out_835,
  output [31:0] io_out_836,
  output [31:0] io_out_837,
  output [31:0] io_out_838,
  output [31:0] io_out_839,
  output [31:0] io_out_840,
  output [31:0] io_out_841,
  output [31:0] io_out_842,
  output [31:0] io_out_843,
  output [31:0] io_out_844,
  output [31:0] io_out_845,
  output [31:0] io_out_846,
  output [31:0] io_out_847,
  output [31:0] io_out_848,
  output [31:0] io_out_849,
  output [31:0] io_out_850,
  output [31:0] io_out_851,
  output [31:0] io_out_852,
  output [31:0] io_out_853,
  output [31:0] io_out_854,
  output [31:0] io_out_855,
  output [31:0] io_out_856,
  output [31:0] io_out_857,
  output [31:0] io_out_858,
  output [31:0] io_out_859,
  output [31:0] io_out_860,
  output [31:0] io_out_861,
  output [31:0] io_out_862,
  output [31:0] io_out_863,
  output [31:0] io_out_864,
  output [31:0] io_out_865,
  output [31:0] io_out_866,
  output [31:0] io_out_867,
  output [31:0] io_out_868,
  output [31:0] io_out_869,
  output [31:0] io_out_870,
  output [31:0] io_out_871,
  output [31:0] io_out_872,
  output [31:0] io_out_873,
  output [31:0] io_out_874,
  output [31:0] io_out_875,
  output [31:0] io_out_876,
  output [31:0] io_out_877,
  output [31:0] io_out_878,
  output [31:0] io_out_879,
  output [31:0] io_out_880,
  output [31:0] io_out_881,
  output [31:0] io_out_882,
  output [31:0] io_out_883,
  output [31:0] io_out_884,
  output [31:0] io_out_885,
  output [31:0] io_out_886,
  output [31:0] io_out_887,
  output [31:0] io_out_888,
  output [31:0] io_out_889,
  output [31:0] io_out_890,
  output [31:0] io_out_891,
  output [31:0] io_out_892,
  output [31:0] io_out_893,
  output [31:0] io_out_894,
  output [31:0] io_out_895,
  output [31:0] io_out_896,
  output [31:0] io_out_897,
  output [31:0] io_out_898,
  output [31:0] io_out_899,
  output [31:0] io_out_900,
  output [31:0] io_out_901,
  output [31:0] io_out_902,
  output [31:0] io_out_903,
  output [31:0] io_out_904,
  output [31:0] io_out_905,
  output [31:0] io_out_906,
  output [31:0] io_out_907,
  output [31:0] io_out_908,
  output [31:0] io_out_909,
  output [31:0] io_out_910,
  output [31:0] io_out_911,
  output [31:0] io_out_912,
  output [31:0] io_out_913,
  output [31:0] io_out_914,
  output [31:0] io_out_915,
  output [31:0] io_out_916,
  output [31:0] io_out_917,
  output [31:0] io_out_918,
  output [31:0] io_out_919,
  output [31:0] io_out_920,
  output [31:0] io_out_921,
  output [31:0] io_out_922,
  output [31:0] io_out_923,
  output [31:0] io_out_924,
  output [31:0] io_out_925,
  output [31:0] io_out_926,
  output [31:0] io_out_927,
  output [31:0] io_out_928,
  output [31:0] io_out_929,
  output [31:0] io_out_930,
  output [31:0] io_out_931,
  output [31:0] io_out_932,
  output [31:0] io_out_933,
  output [31:0] io_out_934,
  output [31:0] io_out_935,
  output [31:0] io_out_936,
  output [31:0] io_out_937,
  output [31:0] io_out_938,
  output [31:0] io_out_939,
  output [31:0] io_out_940,
  output [31:0] io_out_941,
  output [31:0] io_out_942,
  output [31:0] io_out_943,
  output [31:0] io_out_944,
  output [31:0] io_out_945,
  output [31:0] io_out_946,
  output [31:0] io_out_947,
  output [31:0] io_out_948,
  output [31:0] io_out_949,
  output [31:0] io_out_950,
  output [31:0] io_out_951,
  output [31:0] io_out_952,
  output [31:0] io_out_953,
  output [31:0] io_out_954,
  output [31:0] io_out_955,
  output [31:0] io_out_956,
  output [31:0] io_out_957,
  output [31:0] io_out_958,
  output [31:0] io_out_959,
  output [31:0] io_out_960,
  output [31:0] io_out_961,
  output [31:0] io_out_962,
  output [31:0] io_out_963,
  output [31:0] io_out_964,
  output [31:0] io_out_965,
  output [31:0] io_out_966,
  output [31:0] io_out_967,
  output [31:0] io_out_968,
  output [31:0] io_out_969,
  output [31:0] io_out_970,
  output [31:0] io_out_971,
  output [31:0] io_out_972,
  output [31:0] io_out_973,
  output [31:0] io_out_974,
  output [31:0] io_out_975,
  output [31:0] io_out_976,
  output [31:0] io_out_977,
  output [31:0] io_out_978,
  output [31:0] io_out_979,
  output [31:0] io_out_980,
  output [31:0] io_out_981,
  output [31:0] io_out_982,
  output [31:0] io_out_983,
  output [31:0] io_out_984,
  output [31:0] io_out_985,
  output [31:0] io_out_986,
  output [31:0] io_out_987,
  output [31:0] io_out_988,
  output [31:0] io_out_989,
  output [31:0] io_out_990,
  output [31:0] io_out_991,
  output [31:0] io_out_992,
  output [31:0] io_out_993,
  output [31:0] io_out_994,
  output [31:0] io_out_995,
  output [31:0] io_out_996,
  output [31:0] io_out_997,
  output [31:0] io_out_998,
  output [31:0] io_out_999,
  output [31:0] io_out_1000,
  output [31:0] io_out_1001,
  output [31:0] io_out_1002,
  output [31:0] io_out_1003,
  output [31:0] io_out_1004,
  output [31:0] io_out_1005,
  output [31:0] io_out_1006,
  output [31:0] io_out_1007,
  output [31:0] io_out_1008,
  output [31:0] io_out_1009,
  output [31:0] io_out_1010,
  output [31:0] io_out_1011,
  output [31:0] io_out_1012,
  output [31:0] io_out_1013,
  output [31:0] io_out_1014,
  output [31:0] io_out_1015,
  output [31:0] io_out_1016,
  output [31:0] io_out_1017,
  output [31:0] io_out_1018,
  output [31:0] io_out_1019,
  output [31:0] io_out_1020,
  output [31:0] io_out_1021,
  output [31:0] io_out_1022,
  output [31:0] io_out_1023
);
  wire  bc_pe_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_2_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_2_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_2_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_2_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_2_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_2_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_2_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_2_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_2_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_3_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_3_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_3_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_3_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_3_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_3_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_3_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_3_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_3_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_4_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_4_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_4_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_4_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_4_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_4_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_4_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_4_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_4_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_5_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_5_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_5_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_5_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_5_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_5_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_5_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_5_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_5_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_6_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_6_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_6_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_6_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_6_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_6_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_6_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_6_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_6_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_7_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_7_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_7_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_7_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_7_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_7_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_7_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_7_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_7_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_8_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_8_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_8_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_8_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_8_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_8_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_8_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_8_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_8_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_9_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_9_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_9_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_9_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_9_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_9_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_9_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_9_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_9_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_10_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_10_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_10_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_10_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_10_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_10_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_10_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_10_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_10_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_11_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_11_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_11_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_11_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_11_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_11_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_11_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_11_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_11_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_12_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_12_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_12_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_12_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_12_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_12_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_12_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_12_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_12_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_13_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_13_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_13_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_13_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_13_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_13_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_13_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_13_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_13_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_14_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_14_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_14_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_14_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_14_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_14_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_14_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_14_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_14_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_15_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_15_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_15_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_15_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_15_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_15_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_15_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_15_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_15_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_16_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_16_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_16_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_16_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_16_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_16_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_16_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_16_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_16_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_17_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_17_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_17_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_17_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_17_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_17_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_17_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_17_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_17_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_18_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_18_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_18_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_18_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_18_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_18_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_18_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_18_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_18_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_19_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_19_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_19_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_19_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_19_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_19_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_19_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_19_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_19_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_20_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_20_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_20_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_20_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_20_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_20_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_20_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_20_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_20_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_21_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_21_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_21_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_21_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_21_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_21_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_21_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_21_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_21_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_22_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_22_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_22_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_22_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_22_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_22_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_22_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_22_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_22_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_23_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_23_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_23_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_23_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_23_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_23_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_23_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_23_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_23_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_24_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_24_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_24_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_24_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_24_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_24_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_24_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_24_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_24_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_25_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_25_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_25_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_25_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_25_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_25_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_25_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_25_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_25_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_26_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_26_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_26_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_26_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_26_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_26_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_26_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_26_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_26_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_27_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_27_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_27_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_27_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_27_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_27_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_27_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_27_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_27_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_28_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_28_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_28_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_28_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_28_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_28_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_28_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_28_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_28_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_29_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_29_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_29_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_29_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_29_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_29_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_29_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_29_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_29_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_30_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_30_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_30_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_30_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_30_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_30_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_30_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_30_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_30_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_31_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_31_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_31_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_31_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_31_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_31_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_31_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_31_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_31_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_32_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_32_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_32_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_32_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_32_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_32_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_32_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_32_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_32_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_33_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_33_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_33_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_33_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_33_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_33_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_33_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_33_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_33_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_34_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_34_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_34_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_34_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_34_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_34_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_34_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_34_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_34_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_35_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_35_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_35_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_35_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_35_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_35_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_35_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_35_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_35_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_36_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_36_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_36_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_36_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_36_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_36_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_36_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_36_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_36_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_37_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_37_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_37_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_37_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_37_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_37_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_37_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_37_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_37_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_38_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_38_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_38_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_38_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_38_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_38_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_38_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_38_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_38_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_39_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_39_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_39_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_39_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_39_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_39_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_39_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_39_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_39_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_40_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_40_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_40_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_40_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_40_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_40_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_40_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_40_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_40_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_41_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_41_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_41_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_41_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_41_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_41_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_41_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_41_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_41_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_42_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_42_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_42_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_42_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_42_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_42_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_42_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_42_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_42_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_43_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_43_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_43_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_43_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_43_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_43_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_43_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_43_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_43_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_44_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_44_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_44_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_44_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_44_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_44_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_44_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_44_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_44_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_45_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_45_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_45_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_45_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_45_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_45_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_45_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_45_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_45_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_46_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_46_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_46_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_46_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_46_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_46_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_46_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_46_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_46_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_47_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_47_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_47_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_47_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_47_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_47_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_47_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_47_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_47_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_48_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_48_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_48_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_48_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_48_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_48_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_48_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_48_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_48_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_49_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_49_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_49_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_49_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_49_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_49_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_49_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_49_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_49_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_50_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_50_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_50_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_50_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_50_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_50_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_50_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_50_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_50_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_51_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_51_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_51_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_51_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_51_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_51_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_51_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_51_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_51_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_52_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_52_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_52_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_52_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_52_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_52_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_52_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_52_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_52_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_53_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_53_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_53_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_53_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_53_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_53_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_53_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_53_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_53_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_54_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_54_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_54_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_54_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_54_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_54_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_54_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_54_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_54_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_55_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_55_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_55_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_55_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_55_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_55_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_55_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_55_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_55_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_56_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_56_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_56_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_56_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_56_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_56_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_56_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_56_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_56_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_57_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_57_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_57_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_57_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_57_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_57_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_57_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_57_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_57_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_58_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_58_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_58_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_58_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_58_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_58_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_58_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_58_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_58_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_59_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_59_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_59_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_59_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_59_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_59_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_59_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_59_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_59_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_60_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_60_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_60_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_60_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_60_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_60_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_60_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_60_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_60_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_61_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_61_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_61_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_61_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_61_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_61_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_61_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_61_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_61_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_62_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_62_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_62_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_62_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_62_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_62_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_62_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_62_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_62_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_63_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_63_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_63_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_63_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_63_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_63_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_63_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_63_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_63_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_64_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_64_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_64_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_64_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_64_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_64_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_64_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_64_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_64_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_65_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_65_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_65_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_65_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_65_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_65_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_65_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_65_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_65_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_66_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_66_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_66_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_66_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_66_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_66_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_66_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_66_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_66_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_67_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_67_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_67_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_67_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_67_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_67_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_67_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_67_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_67_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_68_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_68_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_68_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_68_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_68_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_68_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_68_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_68_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_68_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_69_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_69_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_69_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_69_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_69_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_69_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_69_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_69_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_69_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_70_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_70_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_70_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_70_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_70_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_70_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_70_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_70_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_70_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_71_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_71_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_71_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_71_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_71_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_71_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_71_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_71_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_71_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_72_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_72_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_72_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_72_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_72_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_72_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_72_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_72_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_72_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_73_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_73_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_73_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_73_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_73_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_73_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_73_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_73_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_73_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_74_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_74_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_74_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_74_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_74_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_74_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_74_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_74_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_74_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_75_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_75_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_75_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_75_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_75_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_75_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_75_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_75_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_75_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_76_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_76_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_76_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_76_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_76_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_76_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_76_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_76_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_76_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_77_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_77_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_77_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_77_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_77_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_77_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_77_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_77_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_77_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_78_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_78_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_78_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_78_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_78_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_78_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_78_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_78_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_78_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_79_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_79_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_79_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_79_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_79_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_79_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_79_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_79_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_79_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_80_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_80_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_80_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_80_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_80_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_80_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_80_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_80_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_80_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_81_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_81_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_81_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_81_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_81_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_81_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_81_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_81_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_81_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_82_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_82_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_82_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_82_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_82_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_82_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_82_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_82_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_82_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_83_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_83_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_83_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_83_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_83_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_83_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_83_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_83_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_83_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_84_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_84_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_84_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_84_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_84_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_84_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_84_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_84_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_84_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_85_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_85_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_85_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_85_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_85_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_85_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_85_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_85_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_85_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_86_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_86_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_86_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_86_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_86_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_86_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_86_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_86_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_86_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_87_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_87_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_87_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_87_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_87_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_87_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_87_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_87_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_87_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_88_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_88_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_88_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_88_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_88_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_88_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_88_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_88_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_88_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_89_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_89_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_89_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_89_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_89_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_89_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_89_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_89_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_89_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_90_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_90_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_90_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_90_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_90_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_90_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_90_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_90_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_90_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_91_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_91_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_91_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_91_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_91_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_91_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_91_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_91_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_91_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_92_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_92_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_92_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_92_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_92_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_92_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_92_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_92_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_92_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_93_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_93_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_93_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_93_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_93_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_93_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_93_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_93_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_93_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_94_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_94_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_94_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_94_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_94_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_94_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_94_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_94_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_94_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_95_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_95_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_95_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_95_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_95_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_95_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_95_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_95_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_95_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_96_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_96_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_96_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_96_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_96_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_96_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_96_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_96_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_96_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_97_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_97_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_97_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_97_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_97_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_97_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_97_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_97_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_97_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_98_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_98_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_98_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_98_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_98_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_98_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_98_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_98_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_98_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_99_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_99_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_99_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_99_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_99_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_99_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_99_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_99_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_99_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_100_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_100_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_100_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_100_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_100_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_100_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_100_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_100_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_100_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_101_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_101_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_101_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_101_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_101_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_101_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_101_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_101_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_101_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_102_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_102_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_102_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_102_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_102_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_102_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_102_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_102_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_102_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_103_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_103_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_103_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_103_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_103_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_103_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_103_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_103_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_103_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_104_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_104_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_104_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_104_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_104_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_104_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_104_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_104_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_104_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_105_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_105_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_105_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_105_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_105_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_105_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_105_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_105_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_105_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_106_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_106_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_106_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_106_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_106_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_106_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_106_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_106_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_106_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_107_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_107_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_107_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_107_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_107_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_107_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_107_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_107_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_107_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_108_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_108_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_108_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_108_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_108_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_108_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_108_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_108_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_108_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_109_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_109_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_109_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_109_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_109_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_109_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_109_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_109_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_109_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_110_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_110_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_110_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_110_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_110_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_110_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_110_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_110_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_110_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_111_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_111_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_111_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_111_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_111_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_111_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_111_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_111_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_111_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_112_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_112_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_112_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_112_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_112_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_112_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_112_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_112_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_112_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_113_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_113_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_113_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_113_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_113_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_113_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_113_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_113_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_113_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_114_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_114_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_114_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_114_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_114_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_114_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_114_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_114_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_114_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_115_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_115_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_115_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_115_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_115_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_115_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_115_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_115_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_115_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_116_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_116_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_116_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_116_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_116_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_116_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_116_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_116_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_116_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_117_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_117_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_117_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_117_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_117_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_117_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_117_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_117_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_117_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_118_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_118_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_118_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_118_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_118_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_118_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_118_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_118_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_118_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_119_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_119_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_119_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_119_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_119_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_119_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_119_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_119_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_119_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_120_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_120_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_120_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_120_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_120_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_120_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_120_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_120_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_120_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_121_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_121_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_121_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_121_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_121_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_121_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_121_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_121_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_121_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_122_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_122_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_122_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_122_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_122_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_122_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_122_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_122_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_122_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_123_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_123_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_123_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_123_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_123_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_123_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_123_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_123_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_123_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_124_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_124_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_124_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_124_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_124_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_124_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_124_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_124_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_124_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_125_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_125_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_125_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_125_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_125_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_125_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_125_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_125_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_125_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_126_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_126_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_126_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_126_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_126_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_126_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_126_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_126_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_126_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_127_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_127_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_127_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_127_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_127_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_127_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_127_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_127_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_127_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_128_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_128_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_128_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_128_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_128_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_128_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_128_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_128_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_128_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_129_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_129_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_129_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_129_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_129_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_129_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_129_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_129_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_129_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_130_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_130_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_130_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_130_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_130_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_130_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_130_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_130_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_130_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_131_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_131_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_131_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_131_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_131_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_131_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_131_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_131_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_131_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_132_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_132_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_132_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_132_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_132_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_132_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_132_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_132_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_132_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_133_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_133_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_133_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_133_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_133_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_133_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_133_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_133_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_133_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_134_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_134_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_134_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_134_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_134_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_134_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_134_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_134_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_134_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_135_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_135_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_135_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_135_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_135_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_135_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_135_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_135_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_135_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_136_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_136_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_136_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_136_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_136_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_136_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_136_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_136_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_136_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_137_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_137_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_137_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_137_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_137_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_137_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_137_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_137_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_137_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_138_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_138_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_138_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_138_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_138_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_138_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_138_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_138_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_138_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_139_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_139_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_139_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_139_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_139_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_139_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_139_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_139_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_139_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_140_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_140_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_140_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_140_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_140_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_140_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_140_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_140_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_140_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_141_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_141_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_141_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_141_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_141_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_141_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_141_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_141_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_141_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_142_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_142_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_142_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_142_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_142_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_142_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_142_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_142_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_142_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_143_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_143_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_143_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_143_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_143_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_143_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_143_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_143_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_143_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_144_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_144_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_144_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_144_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_144_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_144_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_144_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_144_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_144_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_145_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_145_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_145_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_145_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_145_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_145_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_145_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_145_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_145_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_146_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_146_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_146_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_146_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_146_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_146_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_146_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_146_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_146_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_147_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_147_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_147_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_147_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_147_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_147_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_147_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_147_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_147_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_148_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_148_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_148_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_148_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_148_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_148_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_148_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_148_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_148_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_149_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_149_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_149_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_149_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_149_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_149_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_149_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_149_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_149_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_150_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_150_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_150_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_150_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_150_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_150_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_150_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_150_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_150_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_151_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_151_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_151_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_151_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_151_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_151_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_151_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_151_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_151_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_152_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_152_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_152_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_152_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_152_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_152_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_152_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_152_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_152_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_153_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_153_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_153_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_153_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_153_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_153_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_153_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_153_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_153_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_154_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_154_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_154_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_154_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_154_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_154_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_154_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_154_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_154_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_155_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_155_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_155_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_155_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_155_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_155_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_155_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_155_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_155_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_156_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_156_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_156_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_156_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_156_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_156_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_156_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_156_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_156_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_157_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_157_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_157_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_157_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_157_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_157_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_157_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_157_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_157_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_158_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_158_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_158_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_158_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_158_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_158_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_158_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_158_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_158_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_159_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_159_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_159_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_159_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_159_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_159_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_159_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_159_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_159_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_160_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_160_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_160_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_160_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_160_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_160_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_160_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_160_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_160_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_161_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_161_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_161_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_161_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_161_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_161_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_161_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_161_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_161_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_162_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_162_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_162_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_162_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_162_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_162_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_162_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_162_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_162_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_163_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_163_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_163_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_163_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_163_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_163_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_163_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_163_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_163_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_164_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_164_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_164_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_164_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_164_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_164_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_164_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_164_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_164_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_165_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_165_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_165_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_165_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_165_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_165_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_165_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_165_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_165_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_166_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_166_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_166_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_166_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_166_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_166_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_166_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_166_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_166_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_167_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_167_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_167_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_167_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_167_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_167_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_167_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_167_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_167_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_168_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_168_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_168_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_168_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_168_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_168_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_168_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_168_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_168_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_169_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_169_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_169_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_169_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_169_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_169_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_169_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_169_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_169_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_170_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_170_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_170_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_170_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_170_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_170_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_170_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_170_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_170_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_171_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_171_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_171_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_171_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_171_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_171_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_171_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_171_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_171_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_172_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_172_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_172_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_172_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_172_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_172_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_172_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_172_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_172_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_173_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_173_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_173_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_173_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_173_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_173_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_173_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_173_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_173_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_174_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_174_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_174_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_174_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_174_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_174_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_174_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_174_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_174_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_175_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_175_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_175_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_175_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_175_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_175_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_175_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_175_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_175_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_176_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_176_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_176_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_176_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_176_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_176_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_176_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_176_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_176_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_177_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_177_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_177_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_177_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_177_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_177_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_177_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_177_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_177_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_178_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_178_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_178_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_178_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_178_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_178_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_178_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_178_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_178_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_179_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_179_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_179_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_179_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_179_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_179_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_179_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_179_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_179_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_180_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_180_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_180_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_180_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_180_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_180_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_180_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_180_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_180_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_181_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_181_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_181_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_181_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_181_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_181_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_181_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_181_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_181_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_182_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_182_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_182_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_182_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_182_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_182_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_182_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_182_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_182_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_183_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_183_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_183_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_183_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_183_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_183_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_183_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_183_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_183_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_184_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_184_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_184_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_184_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_184_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_184_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_184_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_184_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_184_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_185_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_185_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_185_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_185_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_185_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_185_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_185_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_185_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_185_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_186_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_186_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_186_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_186_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_186_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_186_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_186_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_186_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_186_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_187_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_187_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_187_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_187_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_187_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_187_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_187_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_187_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_187_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_188_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_188_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_188_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_188_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_188_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_188_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_188_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_188_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_188_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_189_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_189_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_189_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_189_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_189_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_189_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_189_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_189_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_189_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_190_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_190_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_190_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_190_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_190_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_190_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_190_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_190_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_190_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_191_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_191_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_191_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_191_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_191_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_191_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_191_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_191_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_191_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_192_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_192_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_192_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_192_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_192_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_192_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_192_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_192_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_192_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_193_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_193_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_193_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_193_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_193_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_193_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_193_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_193_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_193_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_194_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_194_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_194_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_194_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_194_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_194_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_194_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_194_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_194_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_195_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_195_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_195_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_195_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_195_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_195_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_195_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_195_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_195_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_196_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_196_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_196_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_196_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_196_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_196_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_196_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_196_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_196_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_197_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_197_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_197_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_197_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_197_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_197_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_197_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_197_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_197_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_198_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_198_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_198_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_198_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_198_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_198_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_198_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_198_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_198_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_199_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_199_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_199_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_199_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_199_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_199_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_199_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_199_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_199_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_200_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_200_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_200_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_200_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_200_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_200_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_200_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_200_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_200_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_201_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_201_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_201_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_201_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_201_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_201_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_201_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_201_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_201_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_202_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_202_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_202_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_202_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_202_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_202_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_202_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_202_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_202_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_203_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_203_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_203_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_203_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_203_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_203_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_203_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_203_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_203_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_204_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_204_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_204_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_204_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_204_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_204_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_204_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_204_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_204_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_205_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_205_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_205_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_205_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_205_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_205_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_205_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_205_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_205_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_206_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_206_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_206_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_206_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_206_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_206_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_206_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_206_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_206_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_207_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_207_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_207_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_207_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_207_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_207_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_207_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_207_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_207_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_208_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_208_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_208_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_208_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_208_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_208_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_208_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_208_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_208_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_209_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_209_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_209_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_209_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_209_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_209_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_209_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_209_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_209_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_210_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_210_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_210_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_210_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_210_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_210_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_210_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_210_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_210_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_211_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_211_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_211_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_211_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_211_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_211_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_211_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_211_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_211_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_212_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_212_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_212_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_212_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_212_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_212_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_212_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_212_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_212_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_213_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_213_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_213_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_213_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_213_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_213_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_213_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_213_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_213_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_214_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_214_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_214_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_214_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_214_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_214_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_214_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_214_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_214_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_215_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_215_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_215_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_215_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_215_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_215_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_215_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_215_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_215_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_216_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_216_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_216_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_216_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_216_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_216_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_216_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_216_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_216_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_217_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_217_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_217_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_217_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_217_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_217_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_217_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_217_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_217_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_218_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_218_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_218_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_218_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_218_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_218_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_218_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_218_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_218_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_219_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_219_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_219_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_219_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_219_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_219_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_219_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_219_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_219_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_220_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_220_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_220_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_220_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_220_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_220_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_220_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_220_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_220_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_221_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_221_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_221_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_221_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_221_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_221_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_221_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_221_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_221_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_222_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_222_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_222_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_222_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_222_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_222_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_222_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_222_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_222_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_223_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_223_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_223_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_223_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_223_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_223_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_223_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_223_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_223_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_224_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_224_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_224_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_224_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_224_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_224_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_224_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_224_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_224_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_225_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_225_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_225_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_225_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_225_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_225_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_225_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_225_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_225_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_226_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_226_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_226_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_226_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_226_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_226_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_226_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_226_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_226_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_227_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_227_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_227_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_227_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_227_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_227_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_227_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_227_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_227_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_228_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_228_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_228_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_228_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_228_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_228_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_228_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_228_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_228_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_229_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_229_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_229_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_229_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_229_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_229_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_229_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_229_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_229_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_230_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_230_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_230_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_230_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_230_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_230_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_230_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_230_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_230_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_231_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_231_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_231_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_231_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_231_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_231_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_231_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_231_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_231_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_232_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_232_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_232_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_232_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_232_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_232_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_232_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_232_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_232_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_233_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_233_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_233_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_233_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_233_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_233_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_233_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_233_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_233_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_234_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_234_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_234_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_234_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_234_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_234_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_234_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_234_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_234_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_235_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_235_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_235_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_235_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_235_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_235_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_235_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_235_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_235_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_236_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_236_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_236_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_236_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_236_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_236_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_236_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_236_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_236_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_237_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_237_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_237_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_237_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_237_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_237_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_237_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_237_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_237_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_238_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_238_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_238_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_238_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_238_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_238_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_238_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_238_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_238_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_239_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_239_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_239_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_239_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_239_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_239_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_239_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_239_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_239_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_240_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_240_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_240_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_240_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_240_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_240_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_240_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_240_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_240_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_241_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_241_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_241_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_241_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_241_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_241_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_241_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_241_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_241_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_242_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_242_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_242_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_242_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_242_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_242_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_242_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_242_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_242_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_243_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_243_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_243_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_243_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_243_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_243_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_243_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_243_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_243_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_244_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_244_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_244_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_244_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_244_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_244_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_244_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_244_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_244_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_245_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_245_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_245_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_245_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_245_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_245_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_245_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_245_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_245_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_246_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_246_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_246_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_246_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_246_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_246_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_246_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_246_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_246_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_247_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_247_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_247_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_247_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_247_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_247_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_247_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_247_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_247_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_248_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_248_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_248_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_248_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_248_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_248_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_248_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_248_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_248_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_249_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_249_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_249_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_249_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_249_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_249_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_249_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_249_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_249_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_250_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_250_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_250_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_250_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_250_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_250_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_250_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_250_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_250_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_251_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_251_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_251_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_251_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_251_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_251_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_251_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_251_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_251_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_252_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_252_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_252_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_252_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_252_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_252_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_252_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_252_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_252_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_253_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_253_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_253_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_253_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_253_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_253_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_253_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_253_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_253_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_254_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_254_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_254_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_254_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_254_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_254_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_254_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_254_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_254_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_255_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_255_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_255_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_255_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_255_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_255_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_255_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_255_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_255_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_256_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_256_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_256_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_256_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_256_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_256_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_256_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_256_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_256_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_257_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_257_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_257_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_257_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_257_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_257_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_257_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_257_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_257_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_258_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_258_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_258_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_258_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_258_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_258_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_258_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_258_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_258_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_259_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_259_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_259_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_259_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_259_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_259_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_259_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_259_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_259_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_260_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_260_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_260_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_260_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_260_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_260_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_260_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_260_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_260_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_261_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_261_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_261_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_261_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_261_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_261_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_261_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_261_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_261_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_262_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_262_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_262_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_262_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_262_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_262_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_262_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_262_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_262_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_263_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_263_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_263_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_263_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_263_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_263_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_263_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_263_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_263_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_264_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_264_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_264_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_264_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_264_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_264_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_264_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_264_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_264_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_265_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_265_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_265_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_265_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_265_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_265_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_265_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_265_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_265_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_266_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_266_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_266_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_266_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_266_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_266_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_266_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_266_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_266_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_267_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_267_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_267_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_267_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_267_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_267_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_267_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_267_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_267_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_268_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_268_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_268_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_268_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_268_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_268_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_268_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_268_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_268_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_269_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_269_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_269_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_269_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_269_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_269_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_269_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_269_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_269_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_270_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_270_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_270_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_270_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_270_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_270_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_270_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_270_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_270_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_271_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_271_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_271_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_271_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_271_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_271_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_271_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_271_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_271_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_272_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_272_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_272_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_272_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_272_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_272_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_272_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_272_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_272_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_273_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_273_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_273_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_273_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_273_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_273_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_273_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_273_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_273_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_274_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_274_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_274_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_274_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_274_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_274_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_274_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_274_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_274_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_275_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_275_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_275_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_275_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_275_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_275_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_275_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_275_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_275_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_276_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_276_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_276_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_276_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_276_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_276_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_276_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_276_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_276_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_277_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_277_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_277_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_277_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_277_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_277_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_277_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_277_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_277_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_278_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_278_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_278_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_278_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_278_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_278_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_278_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_278_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_278_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_279_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_279_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_279_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_279_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_279_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_279_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_279_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_279_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_279_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_280_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_280_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_280_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_280_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_280_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_280_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_280_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_280_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_280_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_281_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_281_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_281_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_281_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_281_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_281_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_281_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_281_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_281_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_282_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_282_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_282_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_282_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_282_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_282_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_282_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_282_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_282_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_283_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_283_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_283_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_283_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_283_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_283_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_283_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_283_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_283_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_284_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_284_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_284_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_284_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_284_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_284_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_284_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_284_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_284_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_285_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_285_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_285_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_285_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_285_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_285_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_285_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_285_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_285_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_286_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_286_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_286_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_286_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_286_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_286_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_286_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_286_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_286_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_287_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_287_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_287_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_287_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_287_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_287_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_287_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_287_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_287_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_288_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_288_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_288_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_288_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_288_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_288_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_288_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_288_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_288_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_289_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_289_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_289_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_289_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_289_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_289_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_289_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_289_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_289_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_290_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_290_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_290_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_290_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_290_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_290_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_290_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_290_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_290_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_291_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_291_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_291_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_291_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_291_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_291_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_291_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_291_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_291_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_292_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_292_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_292_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_292_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_292_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_292_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_292_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_292_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_292_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_293_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_293_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_293_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_293_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_293_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_293_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_293_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_293_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_293_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_294_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_294_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_294_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_294_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_294_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_294_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_294_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_294_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_294_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_295_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_295_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_295_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_295_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_295_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_295_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_295_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_295_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_295_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_296_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_296_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_296_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_296_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_296_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_296_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_296_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_296_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_296_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_297_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_297_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_297_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_297_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_297_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_297_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_297_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_297_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_297_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_298_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_298_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_298_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_298_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_298_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_298_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_298_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_298_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_298_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_299_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_299_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_299_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_299_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_299_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_299_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_299_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_299_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_299_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_300_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_300_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_300_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_300_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_300_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_300_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_300_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_300_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_300_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_301_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_301_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_301_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_301_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_301_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_301_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_301_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_301_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_301_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_302_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_302_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_302_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_302_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_302_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_302_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_302_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_302_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_302_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_303_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_303_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_303_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_303_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_303_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_303_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_303_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_303_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_303_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_304_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_304_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_304_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_304_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_304_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_304_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_304_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_304_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_304_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_305_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_305_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_305_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_305_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_305_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_305_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_305_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_305_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_305_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_306_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_306_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_306_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_306_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_306_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_306_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_306_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_306_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_306_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_307_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_307_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_307_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_307_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_307_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_307_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_307_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_307_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_307_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_308_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_308_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_308_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_308_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_308_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_308_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_308_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_308_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_308_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_309_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_309_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_309_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_309_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_309_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_309_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_309_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_309_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_309_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_310_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_310_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_310_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_310_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_310_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_310_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_310_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_310_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_310_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_311_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_311_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_311_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_311_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_311_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_311_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_311_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_311_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_311_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_312_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_312_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_312_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_312_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_312_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_312_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_312_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_312_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_312_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_313_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_313_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_313_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_313_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_313_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_313_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_313_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_313_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_313_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_314_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_314_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_314_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_314_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_314_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_314_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_314_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_314_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_314_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_315_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_315_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_315_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_315_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_315_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_315_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_315_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_315_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_315_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_316_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_316_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_316_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_316_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_316_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_316_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_316_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_316_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_316_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_317_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_317_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_317_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_317_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_317_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_317_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_317_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_317_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_317_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_318_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_318_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_318_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_318_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_318_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_318_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_318_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_318_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_318_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_319_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_319_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_319_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_319_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_319_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_319_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_319_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_319_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_319_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_320_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_320_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_320_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_320_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_320_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_320_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_320_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_320_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_320_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_321_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_321_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_321_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_321_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_321_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_321_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_321_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_321_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_321_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_322_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_322_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_322_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_322_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_322_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_322_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_322_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_322_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_322_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_323_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_323_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_323_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_323_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_323_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_323_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_323_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_323_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_323_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_324_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_324_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_324_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_324_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_324_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_324_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_324_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_324_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_324_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_325_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_325_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_325_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_325_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_325_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_325_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_325_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_325_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_325_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_326_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_326_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_326_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_326_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_326_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_326_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_326_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_326_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_326_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_327_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_327_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_327_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_327_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_327_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_327_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_327_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_327_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_327_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_328_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_328_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_328_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_328_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_328_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_328_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_328_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_328_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_328_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_329_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_329_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_329_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_329_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_329_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_329_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_329_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_329_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_329_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_330_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_330_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_330_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_330_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_330_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_330_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_330_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_330_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_330_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_331_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_331_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_331_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_331_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_331_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_331_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_331_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_331_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_331_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_332_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_332_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_332_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_332_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_332_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_332_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_332_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_332_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_332_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_333_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_333_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_333_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_333_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_333_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_333_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_333_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_333_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_333_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_334_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_334_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_334_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_334_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_334_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_334_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_334_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_334_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_334_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_335_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_335_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_335_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_335_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_335_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_335_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_335_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_335_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_335_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_336_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_336_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_336_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_336_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_336_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_336_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_336_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_336_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_336_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_337_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_337_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_337_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_337_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_337_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_337_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_337_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_337_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_337_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_338_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_338_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_338_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_338_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_338_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_338_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_338_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_338_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_338_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_339_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_339_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_339_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_339_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_339_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_339_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_339_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_339_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_339_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_340_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_340_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_340_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_340_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_340_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_340_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_340_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_340_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_340_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_341_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_341_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_341_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_341_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_341_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_341_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_341_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_341_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_341_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_342_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_342_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_342_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_342_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_342_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_342_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_342_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_342_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_342_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_343_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_343_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_343_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_343_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_343_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_343_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_343_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_343_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_343_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_344_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_344_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_344_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_344_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_344_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_344_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_344_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_344_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_344_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_345_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_345_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_345_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_345_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_345_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_345_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_345_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_345_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_345_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_346_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_346_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_346_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_346_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_346_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_346_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_346_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_346_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_346_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_347_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_347_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_347_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_347_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_347_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_347_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_347_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_347_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_347_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_348_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_348_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_348_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_348_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_348_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_348_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_348_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_348_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_348_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_349_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_349_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_349_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_349_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_349_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_349_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_349_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_349_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_349_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_350_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_350_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_350_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_350_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_350_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_350_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_350_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_350_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_350_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_351_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_351_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_351_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_351_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_351_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_351_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_351_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_351_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_351_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_352_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_352_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_352_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_352_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_352_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_352_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_352_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_352_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_352_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_353_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_353_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_353_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_353_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_353_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_353_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_353_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_353_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_353_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_354_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_354_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_354_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_354_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_354_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_354_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_354_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_354_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_354_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_355_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_355_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_355_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_355_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_355_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_355_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_355_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_355_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_355_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_356_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_356_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_356_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_356_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_356_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_356_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_356_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_356_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_356_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_357_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_357_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_357_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_357_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_357_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_357_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_357_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_357_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_357_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_358_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_358_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_358_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_358_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_358_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_358_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_358_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_358_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_358_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_359_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_359_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_359_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_359_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_359_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_359_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_359_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_359_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_359_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_360_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_360_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_360_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_360_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_360_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_360_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_360_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_360_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_360_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_361_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_361_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_361_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_361_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_361_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_361_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_361_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_361_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_361_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_362_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_362_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_362_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_362_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_362_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_362_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_362_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_362_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_362_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_363_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_363_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_363_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_363_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_363_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_363_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_363_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_363_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_363_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_364_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_364_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_364_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_364_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_364_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_364_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_364_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_364_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_364_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_365_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_365_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_365_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_365_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_365_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_365_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_365_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_365_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_365_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_366_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_366_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_366_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_366_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_366_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_366_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_366_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_366_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_366_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_367_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_367_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_367_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_367_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_367_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_367_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_367_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_367_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_367_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_368_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_368_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_368_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_368_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_368_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_368_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_368_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_368_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_368_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_369_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_369_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_369_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_369_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_369_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_369_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_369_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_369_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_369_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_370_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_370_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_370_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_370_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_370_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_370_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_370_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_370_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_370_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_371_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_371_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_371_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_371_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_371_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_371_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_371_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_371_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_371_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_372_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_372_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_372_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_372_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_372_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_372_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_372_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_372_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_372_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_373_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_373_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_373_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_373_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_373_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_373_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_373_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_373_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_373_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_374_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_374_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_374_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_374_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_374_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_374_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_374_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_374_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_374_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_375_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_375_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_375_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_375_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_375_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_375_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_375_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_375_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_375_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_376_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_376_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_376_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_376_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_376_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_376_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_376_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_376_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_376_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_377_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_377_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_377_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_377_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_377_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_377_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_377_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_377_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_377_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_378_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_378_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_378_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_378_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_378_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_378_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_378_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_378_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_378_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_379_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_379_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_379_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_379_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_379_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_379_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_379_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_379_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_379_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_380_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_380_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_380_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_380_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_380_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_380_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_380_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_380_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_380_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_381_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_381_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_381_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_381_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_381_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_381_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_381_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_381_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_381_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_382_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_382_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_382_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_382_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_382_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_382_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_382_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_382_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_382_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_383_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_383_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_383_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_383_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_383_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_383_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_383_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_383_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_383_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_384_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_384_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_384_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_384_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_384_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_384_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_384_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_384_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_384_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_385_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_385_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_385_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_385_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_385_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_385_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_385_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_385_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_385_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_386_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_386_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_386_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_386_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_386_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_386_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_386_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_386_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_386_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_387_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_387_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_387_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_387_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_387_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_387_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_387_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_387_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_387_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_388_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_388_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_388_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_388_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_388_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_388_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_388_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_388_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_388_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_389_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_389_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_389_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_389_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_389_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_389_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_389_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_389_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_389_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_390_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_390_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_390_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_390_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_390_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_390_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_390_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_390_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_390_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_391_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_391_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_391_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_391_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_391_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_391_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_391_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_391_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_391_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_392_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_392_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_392_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_392_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_392_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_392_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_392_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_392_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_392_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_393_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_393_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_393_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_393_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_393_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_393_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_393_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_393_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_393_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_394_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_394_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_394_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_394_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_394_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_394_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_394_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_394_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_394_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_395_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_395_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_395_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_395_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_395_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_395_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_395_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_395_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_395_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_396_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_396_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_396_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_396_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_396_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_396_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_396_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_396_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_396_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_397_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_397_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_397_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_397_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_397_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_397_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_397_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_397_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_397_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_398_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_398_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_398_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_398_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_398_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_398_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_398_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_398_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_398_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_399_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_399_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_399_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_399_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_399_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_399_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_399_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_399_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_399_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_400_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_400_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_400_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_400_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_400_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_400_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_400_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_400_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_400_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_401_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_401_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_401_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_401_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_401_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_401_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_401_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_401_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_401_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_402_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_402_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_402_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_402_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_402_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_402_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_402_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_402_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_402_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_403_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_403_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_403_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_403_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_403_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_403_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_403_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_403_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_403_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_404_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_404_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_404_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_404_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_404_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_404_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_404_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_404_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_404_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_405_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_405_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_405_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_405_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_405_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_405_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_405_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_405_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_405_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_406_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_406_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_406_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_406_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_406_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_406_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_406_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_406_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_406_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_407_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_407_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_407_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_407_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_407_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_407_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_407_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_407_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_407_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_408_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_408_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_408_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_408_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_408_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_408_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_408_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_408_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_408_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_409_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_409_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_409_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_409_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_409_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_409_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_409_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_409_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_409_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_410_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_410_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_410_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_410_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_410_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_410_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_410_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_410_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_410_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_411_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_411_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_411_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_411_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_411_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_411_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_411_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_411_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_411_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_412_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_412_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_412_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_412_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_412_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_412_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_412_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_412_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_412_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_413_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_413_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_413_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_413_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_413_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_413_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_413_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_413_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_413_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_414_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_414_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_414_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_414_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_414_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_414_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_414_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_414_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_414_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_415_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_415_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_415_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_415_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_415_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_415_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_415_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_415_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_415_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_416_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_416_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_416_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_416_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_416_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_416_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_416_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_416_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_416_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_417_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_417_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_417_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_417_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_417_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_417_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_417_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_417_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_417_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_418_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_418_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_418_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_418_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_418_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_418_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_418_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_418_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_418_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_419_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_419_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_419_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_419_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_419_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_419_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_419_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_419_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_419_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_420_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_420_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_420_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_420_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_420_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_420_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_420_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_420_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_420_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_421_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_421_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_421_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_421_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_421_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_421_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_421_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_421_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_421_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_422_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_422_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_422_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_422_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_422_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_422_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_422_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_422_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_422_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_423_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_423_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_423_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_423_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_423_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_423_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_423_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_423_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_423_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_424_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_424_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_424_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_424_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_424_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_424_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_424_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_424_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_424_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_425_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_425_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_425_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_425_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_425_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_425_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_425_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_425_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_425_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_426_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_426_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_426_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_426_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_426_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_426_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_426_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_426_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_426_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_427_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_427_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_427_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_427_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_427_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_427_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_427_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_427_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_427_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_428_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_428_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_428_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_428_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_428_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_428_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_428_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_428_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_428_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_429_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_429_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_429_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_429_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_429_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_429_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_429_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_429_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_429_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_430_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_430_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_430_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_430_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_430_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_430_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_430_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_430_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_430_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_431_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_431_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_431_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_431_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_431_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_431_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_431_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_431_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_431_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_432_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_432_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_432_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_432_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_432_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_432_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_432_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_432_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_432_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_433_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_433_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_433_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_433_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_433_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_433_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_433_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_433_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_433_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_434_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_434_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_434_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_434_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_434_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_434_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_434_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_434_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_434_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_435_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_435_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_435_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_435_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_435_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_435_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_435_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_435_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_435_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_436_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_436_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_436_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_436_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_436_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_436_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_436_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_436_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_436_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_437_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_437_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_437_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_437_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_437_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_437_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_437_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_437_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_437_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_438_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_438_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_438_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_438_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_438_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_438_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_438_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_438_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_438_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_439_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_439_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_439_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_439_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_439_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_439_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_439_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_439_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_439_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_440_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_440_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_440_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_440_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_440_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_440_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_440_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_440_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_440_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_441_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_441_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_441_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_441_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_441_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_441_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_441_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_441_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_441_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_442_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_442_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_442_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_442_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_442_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_442_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_442_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_442_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_442_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_443_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_443_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_443_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_443_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_443_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_443_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_443_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_443_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_443_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_444_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_444_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_444_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_444_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_444_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_444_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_444_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_444_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_444_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_445_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_445_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_445_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_445_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_445_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_445_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_445_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_445_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_445_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_446_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_446_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_446_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_446_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_446_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_446_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_446_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_446_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_446_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_447_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_447_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_447_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_447_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_447_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_447_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_447_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_447_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_447_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_448_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_448_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_448_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_448_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_448_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_448_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_448_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_448_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_448_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_449_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_449_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_449_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_449_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_449_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_449_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_449_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_449_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_449_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_450_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_450_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_450_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_450_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_450_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_450_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_450_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_450_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_450_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_451_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_451_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_451_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_451_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_451_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_451_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_451_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_451_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_451_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_452_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_452_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_452_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_452_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_452_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_452_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_452_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_452_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_452_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_453_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_453_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_453_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_453_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_453_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_453_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_453_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_453_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_453_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_454_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_454_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_454_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_454_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_454_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_454_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_454_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_454_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_454_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_455_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_455_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_455_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_455_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_455_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_455_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_455_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_455_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_455_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_456_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_456_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_456_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_456_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_456_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_456_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_456_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_456_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_456_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_457_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_457_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_457_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_457_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_457_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_457_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_457_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_457_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_457_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_458_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_458_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_458_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_458_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_458_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_458_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_458_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_458_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_458_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_459_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_459_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_459_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_459_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_459_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_459_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_459_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_459_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_459_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_460_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_460_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_460_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_460_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_460_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_460_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_460_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_460_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_460_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_461_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_461_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_461_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_461_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_461_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_461_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_461_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_461_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_461_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_462_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_462_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_462_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_462_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_462_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_462_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_462_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_462_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_462_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_463_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_463_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_463_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_463_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_463_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_463_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_463_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_463_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_463_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_464_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_464_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_464_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_464_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_464_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_464_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_464_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_464_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_464_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_465_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_465_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_465_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_465_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_465_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_465_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_465_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_465_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_465_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_466_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_466_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_466_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_466_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_466_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_466_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_466_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_466_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_466_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_467_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_467_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_467_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_467_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_467_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_467_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_467_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_467_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_467_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_468_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_468_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_468_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_468_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_468_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_468_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_468_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_468_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_468_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_469_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_469_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_469_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_469_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_469_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_469_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_469_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_469_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_469_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_470_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_470_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_470_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_470_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_470_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_470_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_470_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_470_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_470_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_471_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_471_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_471_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_471_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_471_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_471_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_471_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_471_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_471_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_472_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_472_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_472_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_472_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_472_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_472_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_472_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_472_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_472_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_473_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_473_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_473_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_473_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_473_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_473_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_473_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_473_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_473_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_474_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_474_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_474_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_474_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_474_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_474_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_474_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_474_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_474_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_475_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_475_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_475_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_475_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_475_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_475_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_475_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_475_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_475_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_476_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_476_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_476_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_476_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_476_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_476_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_476_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_476_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_476_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_477_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_477_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_477_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_477_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_477_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_477_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_477_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_477_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_477_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_478_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_478_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_478_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_478_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_478_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_478_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_478_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_478_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_478_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_479_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_479_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_479_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_479_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_479_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_479_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_479_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_479_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_479_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_480_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_480_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_480_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_480_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_480_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_480_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_480_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_480_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_480_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_481_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_481_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_481_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_481_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_481_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_481_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_481_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_481_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_481_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_482_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_482_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_482_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_482_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_482_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_482_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_482_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_482_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_482_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_483_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_483_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_483_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_483_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_483_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_483_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_483_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_483_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_483_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_484_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_484_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_484_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_484_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_484_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_484_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_484_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_484_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_484_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_485_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_485_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_485_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_485_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_485_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_485_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_485_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_485_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_485_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_486_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_486_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_486_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_486_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_486_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_486_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_486_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_486_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_486_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_487_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_487_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_487_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_487_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_487_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_487_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_487_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_487_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_487_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_488_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_488_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_488_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_488_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_488_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_488_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_488_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_488_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_488_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_489_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_489_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_489_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_489_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_489_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_489_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_489_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_489_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_489_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_490_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_490_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_490_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_490_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_490_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_490_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_490_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_490_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_490_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_491_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_491_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_491_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_491_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_491_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_491_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_491_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_491_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_491_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_492_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_492_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_492_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_492_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_492_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_492_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_492_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_492_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_492_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_493_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_493_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_493_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_493_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_493_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_493_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_493_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_493_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_493_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_494_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_494_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_494_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_494_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_494_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_494_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_494_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_494_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_494_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_495_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_495_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_495_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_495_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_495_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_495_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_495_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_495_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_495_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_496_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_496_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_496_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_496_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_496_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_496_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_496_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_496_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_496_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_497_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_497_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_497_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_497_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_497_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_497_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_497_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_497_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_497_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_498_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_498_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_498_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_498_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_498_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_498_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_498_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_498_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_498_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_499_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_499_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_499_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_499_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_499_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_499_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_499_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_499_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_499_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_500_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_500_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_500_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_500_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_500_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_500_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_500_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_500_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_500_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_501_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_501_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_501_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_501_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_501_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_501_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_501_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_501_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_501_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_502_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_502_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_502_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_502_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_502_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_502_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_502_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_502_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_502_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_503_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_503_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_503_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_503_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_503_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_503_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_503_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_503_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_503_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_504_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_504_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_504_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_504_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_504_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_504_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_504_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_504_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_504_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_505_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_505_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_505_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_505_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_505_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_505_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_505_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_505_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_505_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_506_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_506_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_506_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_506_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_506_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_506_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_506_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_506_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_506_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_507_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_507_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_507_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_507_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_507_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_507_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_507_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_507_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_507_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_508_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_508_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_508_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_508_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_508_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_508_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_508_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_508_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_508_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_509_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_509_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_509_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_509_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_509_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_509_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_509_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_509_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_509_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_510_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_510_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_510_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_510_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_510_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_510_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_510_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_510_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_510_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_511_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_511_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_511_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_511_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_511_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_511_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_511_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_511_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_511_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_512_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_512_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_512_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_512_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_512_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_512_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_512_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_512_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_512_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_513_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_513_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_513_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_513_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_513_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_513_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_513_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_513_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_513_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_514_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_514_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_514_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_514_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_514_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_514_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_514_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_514_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_514_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_515_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_515_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_515_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_515_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_515_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_515_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_515_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_515_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_515_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_516_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_516_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_516_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_516_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_516_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_516_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_516_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_516_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_516_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_517_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_517_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_517_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_517_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_517_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_517_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_517_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_517_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_517_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_518_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_518_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_518_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_518_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_518_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_518_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_518_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_518_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_518_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_519_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_519_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_519_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_519_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_519_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_519_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_519_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_519_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_519_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_520_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_520_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_520_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_520_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_520_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_520_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_520_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_520_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_520_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_521_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_521_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_521_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_521_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_521_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_521_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_521_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_521_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_521_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_522_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_522_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_522_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_522_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_522_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_522_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_522_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_522_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_522_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_523_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_523_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_523_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_523_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_523_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_523_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_523_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_523_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_523_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_524_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_524_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_524_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_524_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_524_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_524_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_524_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_524_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_524_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_525_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_525_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_525_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_525_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_525_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_525_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_525_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_525_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_525_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_526_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_526_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_526_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_526_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_526_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_526_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_526_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_526_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_526_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_527_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_527_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_527_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_527_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_527_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_527_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_527_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_527_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_527_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_528_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_528_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_528_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_528_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_528_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_528_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_528_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_528_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_528_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_529_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_529_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_529_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_529_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_529_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_529_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_529_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_529_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_529_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_530_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_530_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_530_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_530_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_530_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_530_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_530_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_530_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_530_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_531_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_531_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_531_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_531_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_531_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_531_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_531_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_531_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_531_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_532_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_532_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_532_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_532_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_532_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_532_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_532_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_532_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_532_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_533_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_533_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_533_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_533_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_533_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_533_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_533_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_533_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_533_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_534_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_534_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_534_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_534_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_534_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_534_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_534_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_534_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_534_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_535_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_535_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_535_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_535_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_535_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_535_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_535_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_535_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_535_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_536_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_536_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_536_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_536_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_536_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_536_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_536_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_536_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_536_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_537_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_537_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_537_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_537_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_537_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_537_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_537_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_537_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_537_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_538_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_538_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_538_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_538_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_538_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_538_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_538_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_538_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_538_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_539_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_539_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_539_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_539_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_539_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_539_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_539_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_539_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_539_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_540_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_540_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_540_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_540_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_540_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_540_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_540_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_540_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_540_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_541_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_541_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_541_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_541_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_541_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_541_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_541_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_541_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_541_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_542_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_542_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_542_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_542_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_542_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_542_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_542_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_542_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_542_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_543_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_543_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_543_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_543_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_543_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_543_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_543_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_543_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_543_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_544_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_544_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_544_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_544_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_544_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_544_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_544_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_544_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_544_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_545_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_545_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_545_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_545_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_545_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_545_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_545_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_545_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_545_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_546_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_546_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_546_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_546_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_546_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_546_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_546_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_546_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_546_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_547_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_547_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_547_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_547_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_547_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_547_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_547_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_547_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_547_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_548_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_548_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_548_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_548_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_548_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_548_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_548_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_548_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_548_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_549_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_549_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_549_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_549_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_549_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_549_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_549_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_549_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_549_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_550_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_550_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_550_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_550_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_550_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_550_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_550_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_550_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_550_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_551_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_551_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_551_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_551_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_551_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_551_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_551_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_551_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_551_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_552_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_552_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_552_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_552_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_552_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_552_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_552_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_552_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_552_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_553_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_553_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_553_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_553_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_553_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_553_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_553_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_553_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_553_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_554_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_554_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_554_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_554_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_554_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_554_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_554_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_554_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_554_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_555_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_555_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_555_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_555_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_555_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_555_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_555_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_555_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_555_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_556_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_556_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_556_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_556_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_556_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_556_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_556_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_556_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_556_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_557_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_557_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_557_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_557_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_557_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_557_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_557_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_557_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_557_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_558_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_558_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_558_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_558_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_558_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_558_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_558_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_558_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_558_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_559_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_559_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_559_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_559_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_559_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_559_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_559_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_559_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_559_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_560_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_560_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_560_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_560_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_560_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_560_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_560_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_560_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_560_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_561_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_561_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_561_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_561_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_561_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_561_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_561_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_561_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_561_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_562_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_562_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_562_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_562_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_562_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_562_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_562_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_562_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_562_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_563_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_563_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_563_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_563_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_563_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_563_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_563_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_563_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_563_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_564_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_564_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_564_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_564_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_564_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_564_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_564_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_564_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_564_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_565_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_565_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_565_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_565_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_565_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_565_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_565_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_565_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_565_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_566_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_566_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_566_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_566_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_566_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_566_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_566_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_566_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_566_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_567_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_567_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_567_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_567_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_567_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_567_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_567_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_567_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_567_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_568_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_568_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_568_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_568_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_568_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_568_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_568_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_568_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_568_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_569_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_569_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_569_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_569_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_569_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_569_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_569_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_569_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_569_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_570_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_570_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_570_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_570_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_570_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_570_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_570_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_570_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_570_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_571_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_571_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_571_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_571_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_571_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_571_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_571_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_571_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_571_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_572_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_572_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_572_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_572_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_572_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_572_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_572_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_572_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_572_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_573_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_573_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_573_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_573_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_573_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_573_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_573_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_573_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_573_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_574_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_574_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_574_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_574_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_574_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_574_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_574_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_574_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_574_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_575_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_575_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_575_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_575_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_575_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_575_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_575_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_575_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_575_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_576_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_576_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_576_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_576_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_576_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_576_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_576_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_576_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_576_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_577_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_577_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_577_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_577_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_577_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_577_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_577_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_577_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_577_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_578_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_578_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_578_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_578_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_578_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_578_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_578_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_578_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_578_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_579_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_579_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_579_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_579_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_579_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_579_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_579_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_579_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_579_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_580_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_580_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_580_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_580_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_580_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_580_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_580_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_580_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_580_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_581_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_581_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_581_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_581_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_581_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_581_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_581_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_581_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_581_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_582_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_582_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_582_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_582_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_582_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_582_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_582_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_582_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_582_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_583_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_583_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_583_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_583_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_583_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_583_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_583_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_583_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_583_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_584_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_584_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_584_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_584_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_584_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_584_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_584_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_584_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_584_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_585_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_585_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_585_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_585_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_585_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_585_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_585_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_585_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_585_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_586_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_586_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_586_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_586_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_586_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_586_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_586_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_586_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_586_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_587_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_587_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_587_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_587_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_587_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_587_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_587_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_587_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_587_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_588_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_588_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_588_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_588_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_588_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_588_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_588_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_588_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_588_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_589_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_589_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_589_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_589_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_589_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_589_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_589_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_589_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_589_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_590_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_590_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_590_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_590_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_590_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_590_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_590_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_590_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_590_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_591_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_591_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_591_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_591_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_591_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_591_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_591_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_591_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_591_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_592_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_592_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_592_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_592_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_592_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_592_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_592_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_592_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_592_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_593_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_593_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_593_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_593_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_593_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_593_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_593_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_593_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_593_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_594_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_594_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_594_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_594_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_594_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_594_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_594_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_594_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_594_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_595_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_595_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_595_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_595_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_595_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_595_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_595_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_595_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_595_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_596_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_596_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_596_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_596_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_596_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_596_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_596_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_596_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_596_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_597_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_597_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_597_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_597_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_597_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_597_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_597_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_597_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_597_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_598_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_598_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_598_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_598_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_598_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_598_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_598_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_598_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_598_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_599_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_599_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_599_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_599_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_599_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_599_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_599_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_599_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_599_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_600_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_600_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_600_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_600_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_600_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_600_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_600_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_600_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_600_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_601_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_601_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_601_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_601_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_601_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_601_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_601_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_601_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_601_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_602_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_602_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_602_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_602_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_602_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_602_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_602_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_602_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_602_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_603_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_603_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_603_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_603_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_603_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_603_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_603_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_603_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_603_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_604_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_604_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_604_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_604_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_604_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_604_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_604_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_604_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_604_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_605_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_605_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_605_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_605_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_605_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_605_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_605_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_605_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_605_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_606_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_606_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_606_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_606_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_606_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_606_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_606_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_606_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_606_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_607_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_607_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_607_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_607_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_607_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_607_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_607_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_607_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_607_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_608_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_608_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_608_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_608_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_608_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_608_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_608_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_608_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_608_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_609_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_609_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_609_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_609_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_609_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_609_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_609_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_609_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_609_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_610_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_610_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_610_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_610_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_610_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_610_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_610_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_610_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_610_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_611_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_611_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_611_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_611_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_611_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_611_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_611_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_611_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_611_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_612_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_612_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_612_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_612_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_612_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_612_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_612_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_612_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_612_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_613_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_613_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_613_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_613_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_613_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_613_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_613_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_613_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_613_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_614_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_614_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_614_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_614_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_614_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_614_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_614_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_614_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_614_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_615_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_615_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_615_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_615_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_615_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_615_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_615_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_615_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_615_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_616_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_616_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_616_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_616_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_616_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_616_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_616_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_616_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_616_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_617_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_617_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_617_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_617_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_617_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_617_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_617_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_617_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_617_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_618_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_618_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_618_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_618_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_618_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_618_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_618_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_618_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_618_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_619_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_619_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_619_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_619_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_619_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_619_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_619_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_619_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_619_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_620_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_620_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_620_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_620_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_620_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_620_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_620_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_620_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_620_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_621_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_621_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_621_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_621_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_621_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_621_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_621_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_621_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_621_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_622_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_622_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_622_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_622_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_622_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_622_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_622_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_622_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_622_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_623_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_623_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_623_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_623_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_623_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_623_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_623_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_623_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_623_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_624_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_624_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_624_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_624_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_624_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_624_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_624_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_624_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_624_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_625_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_625_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_625_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_625_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_625_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_625_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_625_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_625_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_625_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_626_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_626_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_626_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_626_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_626_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_626_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_626_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_626_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_626_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_627_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_627_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_627_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_627_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_627_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_627_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_627_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_627_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_627_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_628_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_628_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_628_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_628_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_628_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_628_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_628_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_628_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_628_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_629_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_629_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_629_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_629_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_629_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_629_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_629_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_629_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_629_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_630_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_630_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_630_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_630_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_630_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_630_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_630_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_630_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_630_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_631_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_631_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_631_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_631_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_631_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_631_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_631_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_631_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_631_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_632_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_632_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_632_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_632_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_632_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_632_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_632_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_632_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_632_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_633_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_633_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_633_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_633_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_633_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_633_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_633_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_633_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_633_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_634_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_634_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_634_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_634_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_634_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_634_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_634_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_634_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_634_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_635_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_635_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_635_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_635_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_635_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_635_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_635_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_635_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_635_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_636_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_636_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_636_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_636_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_636_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_636_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_636_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_636_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_636_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_637_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_637_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_637_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_637_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_637_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_637_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_637_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_637_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_637_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_638_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_638_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_638_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_638_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_638_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_638_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_638_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_638_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_638_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_639_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_639_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_639_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_639_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_639_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_639_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_639_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_639_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_639_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_640_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_640_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_640_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_640_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_640_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_640_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_640_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_640_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_640_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_641_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_641_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_641_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_641_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_641_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_641_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_641_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_641_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_641_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_642_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_642_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_642_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_642_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_642_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_642_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_642_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_642_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_642_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_643_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_643_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_643_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_643_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_643_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_643_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_643_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_643_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_643_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_644_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_644_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_644_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_644_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_644_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_644_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_644_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_644_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_644_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_645_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_645_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_645_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_645_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_645_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_645_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_645_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_645_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_645_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_646_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_646_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_646_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_646_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_646_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_646_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_646_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_646_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_646_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_647_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_647_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_647_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_647_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_647_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_647_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_647_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_647_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_647_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_648_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_648_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_648_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_648_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_648_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_648_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_648_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_648_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_648_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_649_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_649_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_649_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_649_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_649_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_649_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_649_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_649_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_649_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_650_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_650_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_650_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_650_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_650_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_650_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_650_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_650_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_650_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_651_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_651_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_651_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_651_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_651_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_651_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_651_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_651_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_651_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_652_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_652_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_652_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_652_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_652_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_652_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_652_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_652_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_652_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_653_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_653_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_653_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_653_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_653_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_653_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_653_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_653_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_653_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_654_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_654_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_654_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_654_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_654_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_654_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_654_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_654_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_654_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_655_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_655_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_655_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_655_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_655_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_655_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_655_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_655_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_655_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_656_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_656_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_656_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_656_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_656_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_656_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_656_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_656_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_656_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_657_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_657_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_657_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_657_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_657_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_657_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_657_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_657_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_657_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_658_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_658_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_658_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_658_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_658_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_658_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_658_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_658_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_658_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_659_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_659_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_659_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_659_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_659_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_659_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_659_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_659_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_659_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_660_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_660_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_660_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_660_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_660_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_660_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_660_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_660_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_660_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_661_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_661_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_661_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_661_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_661_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_661_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_661_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_661_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_661_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_662_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_662_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_662_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_662_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_662_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_662_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_662_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_662_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_662_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_663_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_663_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_663_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_663_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_663_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_663_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_663_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_663_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_663_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_664_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_664_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_664_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_664_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_664_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_664_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_664_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_664_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_664_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_665_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_665_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_665_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_665_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_665_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_665_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_665_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_665_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_665_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_666_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_666_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_666_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_666_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_666_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_666_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_666_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_666_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_666_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_667_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_667_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_667_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_667_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_667_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_667_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_667_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_667_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_667_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_668_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_668_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_668_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_668_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_668_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_668_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_668_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_668_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_668_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_669_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_669_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_669_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_669_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_669_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_669_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_669_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_669_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_669_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_670_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_670_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_670_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_670_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_670_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_670_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_670_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_670_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_670_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_671_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_671_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_671_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_671_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_671_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_671_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_671_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_671_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_671_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_672_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_672_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_672_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_672_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_672_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_672_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_672_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_672_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_672_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_673_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_673_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_673_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_673_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_673_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_673_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_673_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_673_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_673_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_674_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_674_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_674_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_674_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_674_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_674_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_674_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_674_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_674_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_675_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_675_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_675_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_675_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_675_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_675_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_675_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_675_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_675_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_676_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_676_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_676_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_676_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_676_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_676_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_676_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_676_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_676_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_677_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_677_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_677_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_677_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_677_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_677_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_677_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_677_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_677_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_678_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_678_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_678_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_678_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_678_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_678_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_678_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_678_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_678_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_679_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_679_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_679_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_679_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_679_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_679_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_679_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_679_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_679_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_680_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_680_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_680_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_680_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_680_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_680_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_680_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_680_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_680_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_681_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_681_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_681_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_681_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_681_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_681_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_681_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_681_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_681_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_682_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_682_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_682_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_682_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_682_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_682_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_682_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_682_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_682_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_683_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_683_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_683_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_683_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_683_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_683_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_683_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_683_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_683_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_684_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_684_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_684_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_684_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_684_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_684_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_684_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_684_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_684_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_685_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_685_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_685_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_685_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_685_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_685_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_685_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_685_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_685_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_686_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_686_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_686_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_686_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_686_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_686_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_686_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_686_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_686_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_687_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_687_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_687_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_687_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_687_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_687_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_687_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_687_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_687_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_688_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_688_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_688_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_688_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_688_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_688_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_688_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_688_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_688_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_689_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_689_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_689_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_689_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_689_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_689_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_689_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_689_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_689_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_690_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_690_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_690_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_690_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_690_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_690_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_690_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_690_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_690_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_691_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_691_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_691_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_691_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_691_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_691_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_691_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_691_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_691_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_692_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_692_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_692_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_692_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_692_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_692_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_692_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_692_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_692_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_693_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_693_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_693_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_693_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_693_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_693_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_693_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_693_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_693_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_694_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_694_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_694_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_694_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_694_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_694_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_694_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_694_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_694_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_695_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_695_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_695_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_695_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_695_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_695_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_695_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_695_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_695_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_696_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_696_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_696_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_696_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_696_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_696_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_696_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_696_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_696_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_697_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_697_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_697_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_697_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_697_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_697_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_697_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_697_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_697_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_698_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_698_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_698_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_698_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_698_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_698_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_698_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_698_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_698_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_699_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_699_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_699_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_699_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_699_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_699_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_699_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_699_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_699_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_700_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_700_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_700_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_700_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_700_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_700_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_700_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_700_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_700_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_701_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_701_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_701_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_701_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_701_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_701_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_701_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_701_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_701_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_702_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_702_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_702_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_702_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_702_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_702_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_702_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_702_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_702_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_703_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_703_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_703_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_703_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_703_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_703_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_703_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_703_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_703_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_704_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_704_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_704_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_704_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_704_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_704_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_704_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_704_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_704_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_705_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_705_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_705_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_705_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_705_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_705_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_705_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_705_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_705_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_706_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_706_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_706_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_706_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_706_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_706_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_706_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_706_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_706_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_707_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_707_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_707_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_707_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_707_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_707_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_707_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_707_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_707_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_708_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_708_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_708_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_708_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_708_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_708_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_708_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_708_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_708_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_709_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_709_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_709_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_709_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_709_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_709_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_709_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_709_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_709_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_710_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_710_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_710_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_710_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_710_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_710_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_710_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_710_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_710_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_711_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_711_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_711_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_711_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_711_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_711_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_711_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_711_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_711_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_712_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_712_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_712_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_712_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_712_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_712_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_712_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_712_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_712_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_713_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_713_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_713_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_713_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_713_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_713_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_713_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_713_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_713_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_714_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_714_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_714_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_714_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_714_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_714_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_714_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_714_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_714_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_715_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_715_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_715_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_715_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_715_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_715_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_715_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_715_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_715_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_716_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_716_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_716_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_716_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_716_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_716_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_716_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_716_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_716_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_717_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_717_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_717_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_717_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_717_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_717_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_717_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_717_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_717_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_718_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_718_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_718_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_718_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_718_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_718_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_718_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_718_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_718_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_719_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_719_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_719_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_719_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_719_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_719_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_719_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_719_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_719_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_720_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_720_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_720_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_720_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_720_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_720_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_720_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_720_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_720_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_721_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_721_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_721_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_721_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_721_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_721_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_721_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_721_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_721_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_722_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_722_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_722_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_722_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_722_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_722_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_722_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_722_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_722_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_723_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_723_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_723_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_723_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_723_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_723_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_723_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_723_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_723_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_724_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_724_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_724_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_724_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_724_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_724_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_724_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_724_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_724_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_725_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_725_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_725_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_725_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_725_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_725_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_725_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_725_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_725_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_726_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_726_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_726_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_726_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_726_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_726_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_726_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_726_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_726_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_727_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_727_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_727_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_727_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_727_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_727_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_727_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_727_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_727_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_728_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_728_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_728_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_728_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_728_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_728_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_728_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_728_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_728_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_729_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_729_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_729_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_729_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_729_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_729_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_729_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_729_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_729_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_730_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_730_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_730_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_730_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_730_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_730_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_730_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_730_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_730_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_731_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_731_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_731_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_731_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_731_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_731_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_731_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_731_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_731_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_732_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_732_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_732_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_732_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_732_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_732_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_732_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_732_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_732_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_733_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_733_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_733_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_733_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_733_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_733_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_733_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_733_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_733_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_734_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_734_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_734_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_734_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_734_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_734_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_734_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_734_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_734_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_735_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_735_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_735_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_735_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_735_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_735_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_735_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_735_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_735_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_736_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_736_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_736_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_736_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_736_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_736_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_736_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_736_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_736_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_737_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_737_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_737_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_737_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_737_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_737_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_737_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_737_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_737_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_738_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_738_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_738_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_738_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_738_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_738_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_738_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_738_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_738_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_739_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_739_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_739_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_739_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_739_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_739_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_739_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_739_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_739_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_740_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_740_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_740_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_740_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_740_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_740_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_740_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_740_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_740_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_741_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_741_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_741_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_741_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_741_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_741_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_741_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_741_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_741_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_742_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_742_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_742_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_742_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_742_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_742_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_742_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_742_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_742_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_743_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_743_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_743_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_743_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_743_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_743_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_743_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_743_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_743_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_744_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_744_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_744_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_744_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_744_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_744_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_744_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_744_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_744_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_745_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_745_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_745_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_745_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_745_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_745_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_745_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_745_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_745_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_746_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_746_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_746_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_746_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_746_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_746_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_746_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_746_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_746_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_747_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_747_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_747_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_747_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_747_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_747_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_747_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_747_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_747_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_748_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_748_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_748_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_748_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_748_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_748_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_748_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_748_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_748_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_749_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_749_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_749_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_749_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_749_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_749_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_749_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_749_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_749_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_750_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_750_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_750_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_750_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_750_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_750_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_750_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_750_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_750_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_751_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_751_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_751_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_751_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_751_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_751_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_751_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_751_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_751_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_752_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_752_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_752_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_752_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_752_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_752_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_752_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_752_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_752_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_753_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_753_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_753_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_753_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_753_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_753_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_753_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_753_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_753_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_754_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_754_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_754_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_754_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_754_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_754_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_754_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_754_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_754_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_755_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_755_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_755_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_755_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_755_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_755_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_755_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_755_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_755_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_756_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_756_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_756_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_756_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_756_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_756_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_756_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_756_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_756_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_757_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_757_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_757_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_757_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_757_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_757_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_757_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_757_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_757_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_758_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_758_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_758_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_758_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_758_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_758_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_758_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_758_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_758_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_759_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_759_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_759_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_759_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_759_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_759_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_759_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_759_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_759_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_760_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_760_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_760_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_760_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_760_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_760_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_760_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_760_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_760_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_761_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_761_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_761_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_761_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_761_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_761_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_761_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_761_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_761_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_762_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_762_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_762_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_762_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_762_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_762_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_762_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_762_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_762_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_763_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_763_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_763_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_763_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_763_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_763_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_763_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_763_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_763_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_764_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_764_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_764_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_764_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_764_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_764_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_764_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_764_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_764_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_765_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_765_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_765_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_765_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_765_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_765_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_765_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_765_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_765_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_766_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_766_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_766_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_766_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_766_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_766_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_766_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_766_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_766_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_767_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_767_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_767_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_767_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_767_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_767_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_767_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_767_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_767_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_768_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_768_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_768_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_768_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_768_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_768_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_768_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_768_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_768_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_769_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_769_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_769_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_769_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_769_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_769_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_769_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_769_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_769_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_770_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_770_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_770_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_770_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_770_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_770_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_770_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_770_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_770_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_771_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_771_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_771_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_771_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_771_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_771_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_771_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_771_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_771_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_772_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_772_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_772_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_772_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_772_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_772_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_772_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_772_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_772_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_773_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_773_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_773_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_773_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_773_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_773_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_773_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_773_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_773_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_774_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_774_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_774_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_774_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_774_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_774_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_774_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_774_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_774_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_775_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_775_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_775_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_775_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_775_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_775_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_775_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_775_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_775_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_776_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_776_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_776_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_776_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_776_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_776_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_776_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_776_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_776_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_777_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_777_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_777_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_777_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_777_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_777_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_777_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_777_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_777_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_778_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_778_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_778_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_778_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_778_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_778_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_778_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_778_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_778_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_779_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_779_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_779_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_779_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_779_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_779_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_779_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_779_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_779_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_780_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_780_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_780_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_780_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_780_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_780_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_780_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_780_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_780_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_781_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_781_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_781_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_781_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_781_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_781_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_781_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_781_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_781_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_782_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_782_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_782_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_782_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_782_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_782_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_782_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_782_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_782_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_783_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_783_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_783_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_783_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_783_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_783_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_783_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_783_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_783_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_784_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_784_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_784_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_784_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_784_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_784_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_784_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_784_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_784_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_785_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_785_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_785_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_785_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_785_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_785_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_785_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_785_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_785_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_786_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_786_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_786_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_786_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_786_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_786_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_786_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_786_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_786_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_787_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_787_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_787_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_787_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_787_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_787_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_787_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_787_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_787_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_788_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_788_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_788_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_788_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_788_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_788_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_788_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_788_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_788_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_789_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_789_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_789_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_789_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_789_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_789_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_789_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_789_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_789_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_790_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_790_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_790_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_790_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_790_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_790_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_790_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_790_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_790_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_791_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_791_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_791_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_791_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_791_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_791_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_791_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_791_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_791_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_792_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_792_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_792_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_792_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_792_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_792_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_792_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_792_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_792_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_793_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_793_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_793_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_793_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_793_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_793_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_793_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_793_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_793_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_794_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_794_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_794_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_794_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_794_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_794_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_794_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_794_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_794_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_795_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_795_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_795_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_795_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_795_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_795_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_795_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_795_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_795_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_796_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_796_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_796_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_796_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_796_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_796_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_796_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_796_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_796_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_797_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_797_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_797_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_797_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_797_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_797_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_797_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_797_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_797_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_798_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_798_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_798_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_798_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_798_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_798_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_798_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_798_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_798_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_799_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_799_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_799_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_799_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_799_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_799_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_799_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_799_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_799_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_800_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_800_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_800_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_800_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_800_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_800_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_800_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_800_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_800_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_801_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_801_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_801_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_801_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_801_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_801_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_801_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_801_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_801_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_802_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_802_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_802_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_802_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_802_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_802_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_802_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_802_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_802_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_803_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_803_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_803_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_803_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_803_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_803_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_803_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_803_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_803_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_804_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_804_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_804_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_804_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_804_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_804_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_804_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_804_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_804_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_805_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_805_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_805_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_805_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_805_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_805_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_805_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_805_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_805_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_806_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_806_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_806_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_806_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_806_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_806_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_806_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_806_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_806_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_807_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_807_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_807_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_807_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_807_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_807_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_807_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_807_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_807_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_808_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_808_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_808_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_808_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_808_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_808_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_808_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_808_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_808_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_809_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_809_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_809_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_809_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_809_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_809_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_809_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_809_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_809_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_810_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_810_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_810_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_810_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_810_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_810_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_810_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_810_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_810_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_811_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_811_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_811_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_811_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_811_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_811_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_811_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_811_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_811_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_812_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_812_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_812_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_812_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_812_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_812_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_812_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_812_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_812_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_813_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_813_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_813_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_813_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_813_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_813_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_813_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_813_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_813_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_814_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_814_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_814_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_814_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_814_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_814_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_814_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_814_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_814_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_815_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_815_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_815_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_815_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_815_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_815_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_815_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_815_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_815_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_816_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_816_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_816_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_816_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_816_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_816_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_816_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_816_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_816_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_817_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_817_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_817_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_817_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_817_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_817_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_817_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_817_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_817_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_818_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_818_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_818_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_818_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_818_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_818_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_818_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_818_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_818_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_819_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_819_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_819_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_819_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_819_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_819_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_819_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_819_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_819_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_820_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_820_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_820_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_820_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_820_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_820_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_820_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_820_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_820_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_821_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_821_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_821_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_821_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_821_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_821_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_821_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_821_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_821_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_822_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_822_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_822_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_822_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_822_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_822_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_822_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_822_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_822_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_823_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_823_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_823_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_823_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_823_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_823_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_823_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_823_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_823_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_824_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_824_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_824_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_824_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_824_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_824_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_824_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_824_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_824_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_825_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_825_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_825_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_825_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_825_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_825_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_825_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_825_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_825_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_826_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_826_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_826_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_826_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_826_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_826_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_826_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_826_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_826_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_827_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_827_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_827_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_827_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_827_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_827_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_827_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_827_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_827_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_828_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_828_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_828_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_828_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_828_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_828_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_828_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_828_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_828_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_829_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_829_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_829_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_829_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_829_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_829_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_829_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_829_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_829_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_830_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_830_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_830_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_830_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_830_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_830_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_830_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_830_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_830_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_831_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_831_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_831_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_831_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_831_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_831_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_831_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_831_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_831_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_832_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_832_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_832_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_832_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_832_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_832_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_832_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_832_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_832_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_833_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_833_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_833_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_833_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_833_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_833_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_833_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_833_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_833_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_834_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_834_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_834_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_834_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_834_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_834_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_834_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_834_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_834_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_835_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_835_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_835_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_835_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_835_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_835_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_835_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_835_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_835_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_836_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_836_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_836_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_836_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_836_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_836_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_836_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_836_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_836_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_837_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_837_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_837_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_837_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_837_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_837_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_837_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_837_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_837_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_838_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_838_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_838_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_838_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_838_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_838_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_838_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_838_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_838_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_839_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_839_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_839_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_839_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_839_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_839_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_839_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_839_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_839_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_840_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_840_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_840_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_840_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_840_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_840_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_840_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_840_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_840_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_841_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_841_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_841_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_841_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_841_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_841_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_841_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_841_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_841_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_842_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_842_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_842_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_842_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_842_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_842_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_842_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_842_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_842_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_843_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_843_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_843_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_843_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_843_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_843_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_843_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_843_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_843_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_844_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_844_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_844_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_844_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_844_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_844_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_844_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_844_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_844_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_845_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_845_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_845_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_845_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_845_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_845_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_845_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_845_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_845_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_846_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_846_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_846_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_846_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_846_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_846_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_846_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_846_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_846_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_847_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_847_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_847_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_847_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_847_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_847_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_847_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_847_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_847_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_848_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_848_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_848_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_848_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_848_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_848_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_848_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_848_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_848_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_849_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_849_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_849_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_849_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_849_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_849_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_849_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_849_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_849_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_850_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_850_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_850_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_850_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_850_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_850_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_850_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_850_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_850_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_851_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_851_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_851_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_851_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_851_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_851_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_851_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_851_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_851_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_852_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_852_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_852_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_852_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_852_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_852_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_852_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_852_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_852_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_853_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_853_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_853_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_853_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_853_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_853_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_853_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_853_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_853_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_854_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_854_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_854_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_854_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_854_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_854_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_854_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_854_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_854_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_855_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_855_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_855_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_855_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_855_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_855_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_855_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_855_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_855_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_856_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_856_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_856_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_856_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_856_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_856_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_856_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_856_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_856_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_857_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_857_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_857_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_857_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_857_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_857_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_857_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_857_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_857_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_858_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_858_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_858_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_858_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_858_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_858_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_858_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_858_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_858_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_859_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_859_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_859_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_859_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_859_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_859_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_859_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_859_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_859_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_860_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_860_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_860_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_860_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_860_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_860_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_860_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_860_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_860_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_861_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_861_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_861_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_861_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_861_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_861_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_861_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_861_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_861_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_862_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_862_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_862_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_862_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_862_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_862_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_862_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_862_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_862_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_863_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_863_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_863_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_863_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_863_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_863_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_863_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_863_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_863_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_864_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_864_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_864_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_864_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_864_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_864_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_864_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_864_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_864_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_865_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_865_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_865_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_865_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_865_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_865_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_865_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_865_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_865_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_866_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_866_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_866_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_866_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_866_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_866_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_866_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_866_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_866_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_867_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_867_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_867_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_867_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_867_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_867_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_867_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_867_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_867_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_868_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_868_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_868_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_868_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_868_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_868_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_868_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_868_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_868_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_869_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_869_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_869_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_869_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_869_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_869_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_869_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_869_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_869_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_870_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_870_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_870_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_870_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_870_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_870_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_870_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_870_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_870_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_871_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_871_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_871_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_871_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_871_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_871_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_871_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_871_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_871_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_872_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_872_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_872_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_872_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_872_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_872_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_872_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_872_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_872_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_873_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_873_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_873_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_873_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_873_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_873_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_873_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_873_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_873_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_874_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_874_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_874_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_874_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_874_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_874_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_874_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_874_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_874_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_875_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_875_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_875_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_875_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_875_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_875_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_875_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_875_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_875_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_876_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_876_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_876_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_876_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_876_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_876_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_876_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_876_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_876_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_877_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_877_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_877_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_877_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_877_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_877_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_877_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_877_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_877_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_878_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_878_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_878_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_878_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_878_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_878_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_878_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_878_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_878_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_879_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_879_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_879_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_879_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_879_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_879_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_879_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_879_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_879_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_880_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_880_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_880_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_880_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_880_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_880_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_880_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_880_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_880_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_881_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_881_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_881_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_881_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_881_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_881_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_881_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_881_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_881_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_882_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_882_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_882_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_882_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_882_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_882_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_882_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_882_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_882_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_883_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_883_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_883_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_883_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_883_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_883_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_883_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_883_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_883_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_884_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_884_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_884_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_884_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_884_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_884_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_884_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_884_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_884_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_885_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_885_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_885_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_885_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_885_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_885_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_885_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_885_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_885_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_886_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_886_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_886_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_886_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_886_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_886_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_886_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_886_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_886_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_887_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_887_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_887_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_887_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_887_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_887_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_887_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_887_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_887_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_888_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_888_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_888_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_888_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_888_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_888_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_888_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_888_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_888_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_889_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_889_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_889_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_889_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_889_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_889_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_889_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_889_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_889_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_890_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_890_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_890_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_890_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_890_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_890_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_890_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_890_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_890_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_891_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_891_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_891_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_891_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_891_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_891_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_891_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_891_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_891_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_892_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_892_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_892_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_892_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_892_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_892_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_892_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_892_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_892_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_893_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_893_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_893_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_893_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_893_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_893_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_893_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_893_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_893_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_894_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_894_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_894_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_894_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_894_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_894_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_894_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_894_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_894_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_895_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_895_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_895_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_895_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_895_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_895_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_895_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_895_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_895_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_896_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_896_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_896_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_896_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_896_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_896_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_896_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_896_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_896_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_897_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_897_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_897_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_897_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_897_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_897_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_897_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_897_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_897_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_898_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_898_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_898_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_898_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_898_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_898_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_898_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_898_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_898_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_899_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_899_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_899_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_899_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_899_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_899_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_899_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_899_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_899_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_900_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_900_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_900_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_900_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_900_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_900_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_900_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_900_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_900_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_901_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_901_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_901_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_901_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_901_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_901_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_901_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_901_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_901_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_902_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_902_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_902_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_902_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_902_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_902_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_902_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_902_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_902_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_903_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_903_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_903_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_903_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_903_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_903_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_903_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_903_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_903_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_904_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_904_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_904_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_904_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_904_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_904_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_904_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_904_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_904_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_905_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_905_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_905_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_905_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_905_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_905_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_905_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_905_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_905_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_906_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_906_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_906_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_906_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_906_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_906_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_906_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_906_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_906_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_907_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_907_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_907_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_907_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_907_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_907_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_907_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_907_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_907_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_908_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_908_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_908_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_908_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_908_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_908_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_908_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_908_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_908_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_909_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_909_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_909_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_909_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_909_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_909_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_909_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_909_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_909_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_910_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_910_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_910_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_910_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_910_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_910_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_910_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_910_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_910_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_911_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_911_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_911_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_911_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_911_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_911_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_911_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_911_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_911_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_912_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_912_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_912_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_912_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_912_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_912_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_912_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_912_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_912_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_913_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_913_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_913_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_913_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_913_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_913_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_913_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_913_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_913_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_914_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_914_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_914_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_914_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_914_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_914_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_914_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_914_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_914_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_915_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_915_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_915_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_915_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_915_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_915_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_915_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_915_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_915_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_916_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_916_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_916_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_916_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_916_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_916_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_916_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_916_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_916_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_917_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_917_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_917_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_917_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_917_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_917_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_917_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_917_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_917_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_918_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_918_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_918_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_918_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_918_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_918_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_918_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_918_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_918_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_919_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_919_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_919_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_919_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_919_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_919_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_919_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_919_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_919_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_920_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_920_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_920_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_920_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_920_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_920_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_920_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_920_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_920_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_921_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_921_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_921_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_921_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_921_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_921_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_921_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_921_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_921_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_922_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_922_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_922_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_922_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_922_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_922_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_922_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_922_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_922_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_923_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_923_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_923_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_923_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_923_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_923_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_923_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_923_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_923_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_924_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_924_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_924_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_924_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_924_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_924_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_924_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_924_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_924_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_925_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_925_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_925_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_925_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_925_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_925_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_925_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_925_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_925_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_926_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_926_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_926_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_926_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_926_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_926_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_926_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_926_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_926_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_927_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_927_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_927_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_927_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_927_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_927_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_927_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_927_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_927_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_928_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_928_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_928_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_928_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_928_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_928_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_928_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_928_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_928_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_929_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_929_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_929_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_929_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_929_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_929_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_929_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_929_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_929_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_930_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_930_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_930_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_930_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_930_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_930_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_930_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_930_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_930_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_931_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_931_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_931_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_931_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_931_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_931_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_931_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_931_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_931_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_932_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_932_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_932_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_932_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_932_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_932_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_932_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_932_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_932_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_933_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_933_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_933_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_933_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_933_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_933_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_933_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_933_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_933_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_934_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_934_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_934_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_934_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_934_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_934_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_934_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_934_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_934_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_935_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_935_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_935_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_935_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_935_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_935_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_935_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_935_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_935_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_936_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_936_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_936_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_936_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_936_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_936_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_936_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_936_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_936_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_937_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_937_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_937_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_937_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_937_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_937_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_937_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_937_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_937_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_938_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_938_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_938_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_938_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_938_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_938_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_938_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_938_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_938_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_939_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_939_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_939_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_939_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_939_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_939_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_939_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_939_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_939_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_940_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_940_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_940_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_940_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_940_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_940_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_940_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_940_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_940_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_941_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_941_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_941_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_941_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_941_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_941_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_941_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_941_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_941_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_942_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_942_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_942_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_942_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_942_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_942_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_942_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_942_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_942_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_943_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_943_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_943_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_943_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_943_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_943_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_943_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_943_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_943_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_944_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_944_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_944_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_944_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_944_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_944_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_944_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_944_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_944_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_945_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_945_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_945_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_945_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_945_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_945_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_945_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_945_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_945_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_946_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_946_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_946_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_946_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_946_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_946_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_946_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_946_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_946_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_947_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_947_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_947_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_947_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_947_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_947_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_947_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_947_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_947_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_948_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_948_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_948_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_948_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_948_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_948_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_948_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_948_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_948_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_949_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_949_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_949_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_949_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_949_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_949_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_949_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_949_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_949_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_950_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_950_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_950_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_950_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_950_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_950_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_950_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_950_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_950_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_951_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_951_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_951_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_951_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_951_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_951_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_951_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_951_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_951_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_952_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_952_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_952_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_952_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_952_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_952_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_952_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_952_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_952_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_953_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_953_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_953_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_953_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_953_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_953_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_953_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_953_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_953_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_954_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_954_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_954_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_954_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_954_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_954_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_954_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_954_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_954_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_955_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_955_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_955_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_955_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_955_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_955_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_955_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_955_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_955_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_956_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_956_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_956_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_956_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_956_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_956_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_956_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_956_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_956_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_957_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_957_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_957_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_957_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_957_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_957_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_957_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_957_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_957_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_958_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_958_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_958_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_958_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_958_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_958_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_958_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_958_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_958_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_959_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_959_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_959_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_959_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_959_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_959_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_959_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_959_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_959_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_960_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_960_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_960_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_960_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_960_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_960_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_960_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_960_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_960_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_961_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_961_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_961_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_961_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_961_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_961_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_961_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_961_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_961_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_962_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_962_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_962_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_962_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_962_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_962_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_962_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_962_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_962_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_963_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_963_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_963_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_963_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_963_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_963_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_963_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_963_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_963_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_964_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_964_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_964_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_964_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_964_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_964_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_964_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_964_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_964_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_965_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_965_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_965_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_965_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_965_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_965_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_965_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_965_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_965_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_966_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_966_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_966_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_966_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_966_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_966_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_966_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_966_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_966_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_967_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_967_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_967_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_967_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_967_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_967_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_967_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_967_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_967_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_968_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_968_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_968_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_968_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_968_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_968_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_968_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_968_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_968_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_969_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_969_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_969_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_969_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_969_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_969_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_969_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_969_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_969_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_970_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_970_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_970_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_970_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_970_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_970_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_970_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_970_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_970_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_971_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_971_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_971_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_971_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_971_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_971_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_971_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_971_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_971_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_972_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_972_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_972_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_972_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_972_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_972_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_972_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_972_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_972_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_973_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_973_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_973_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_973_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_973_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_973_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_973_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_973_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_973_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_974_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_974_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_974_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_974_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_974_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_974_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_974_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_974_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_974_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_975_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_975_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_975_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_975_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_975_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_975_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_975_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_975_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_975_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_976_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_976_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_976_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_976_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_976_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_976_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_976_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_976_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_976_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_977_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_977_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_977_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_977_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_977_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_977_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_977_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_977_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_977_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_978_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_978_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_978_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_978_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_978_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_978_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_978_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_978_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_978_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_979_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_979_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_979_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_979_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_979_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_979_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_979_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_979_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_979_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_980_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_980_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_980_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_980_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_980_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_980_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_980_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_980_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_980_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_981_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_981_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_981_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_981_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_981_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_981_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_981_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_981_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_981_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_982_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_982_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_982_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_982_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_982_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_982_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_982_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_982_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_982_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_983_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_983_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_983_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_983_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_983_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_983_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_983_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_983_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_983_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_984_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_984_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_984_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_984_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_984_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_984_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_984_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_984_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_984_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_985_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_985_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_985_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_985_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_985_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_985_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_985_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_985_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_985_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_986_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_986_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_986_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_986_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_986_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_986_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_986_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_986_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_986_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_987_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_987_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_987_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_987_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_987_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_987_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_987_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_987_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_987_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_988_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_988_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_988_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_988_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_988_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_988_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_988_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_988_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_988_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_989_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_989_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_989_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_989_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_989_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_989_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_989_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_989_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_989_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_990_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_990_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_990_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_990_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_990_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_990_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_990_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_990_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_990_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_991_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_991_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_991_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_991_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_991_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_991_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_991_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_991_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_991_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_992_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_992_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_992_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_992_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_992_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_992_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_992_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_992_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_992_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_993_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_993_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_993_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_993_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_993_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_993_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_993_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_993_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_993_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_994_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_994_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_994_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_994_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_994_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_994_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_994_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_994_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_994_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_995_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_995_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_995_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_995_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_995_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_995_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_995_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_995_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_995_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_996_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_996_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_996_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_996_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_996_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_996_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_996_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_996_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_996_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_997_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_997_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_997_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_997_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_997_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_997_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_997_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_997_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_997_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_998_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_998_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_998_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_998_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_998_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_998_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_998_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_998_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_998_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_999_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_999_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_999_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_999_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_999_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_999_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_999_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_999_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_999_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1000_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1000_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1000_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1000_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1000_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1000_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1000_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1000_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1000_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1001_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1001_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1001_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1001_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1001_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1001_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1001_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1001_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1001_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1002_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1002_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1002_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1002_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1002_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1002_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1002_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1002_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1002_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1003_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1003_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1003_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1003_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1003_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1003_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1003_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1003_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1003_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1004_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1004_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1004_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1004_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1004_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1004_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1004_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1004_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1004_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1005_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1005_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1005_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1005_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1005_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1005_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1005_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1005_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1005_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1006_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1006_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1006_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1006_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1006_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1006_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1006_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1006_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1006_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1007_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1007_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1007_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1007_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1007_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1007_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1007_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1007_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1007_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1008_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1008_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1008_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1008_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1008_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1008_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1008_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1008_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1008_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1009_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1009_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1009_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1009_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1009_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1009_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1009_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1009_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1009_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1010_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1010_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1010_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1010_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1010_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1010_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1010_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1010_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1010_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1011_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1011_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1011_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1011_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1011_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1011_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1011_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1011_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1011_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1012_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1012_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1012_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1012_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1012_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1012_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1012_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1012_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1012_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1013_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1013_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1013_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1013_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1013_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1013_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1013_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1013_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1013_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1014_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1014_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1014_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1014_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1014_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1014_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1014_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1014_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1014_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1015_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1015_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1015_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1015_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1015_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1015_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1015_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1015_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1015_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1016_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1016_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1016_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1016_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1016_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1016_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1016_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1016_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1016_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1017_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1017_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1017_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1017_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1017_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1017_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1017_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1017_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1017_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1018_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1018_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1018_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1018_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1018_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1018_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1018_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1018_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1018_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1019_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1019_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1019_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1019_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1019_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1019_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1019_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1019_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1019_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1020_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1020_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1020_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1020_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1020_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1020_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1020_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1020_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1020_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1021_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1021_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1021_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1021_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1021_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1021_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1021_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1021_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1021_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1022_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1022_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1022_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1022_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1022_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1022_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1022_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1022_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1022_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1023_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1023_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1023_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1023_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1023_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1023_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1023_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1023_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1023_io_res_out; // @[bc_mmul.scala 23:11]
  bc_pe bc_pe ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_clock),
    .reset(bc_pe_reset),
    .io_ho_input(bc_pe_io_ho_input),
    .io_ve_input(bc_pe_io_ve_input),
    .io_input_valid(bc_pe_io_input_valid),
    .io_iormac(bc_pe_io_iormac),
    .io_ve_out(bc_pe_io_ve_out),
    .io_ho_out(bc_pe_io_ho_out),
    .io_res_out(bc_pe_io_res_out)
  );
  bc_pe bc_pe_1 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1_clock),
    .reset(bc_pe_1_reset),
    .io_ho_input(bc_pe_1_io_ho_input),
    .io_ve_input(bc_pe_1_io_ve_input),
    .io_input_valid(bc_pe_1_io_input_valid),
    .io_iormac(bc_pe_1_io_iormac),
    .io_ve_out(bc_pe_1_io_ve_out),
    .io_ho_out(bc_pe_1_io_ho_out),
    .io_res_out(bc_pe_1_io_res_out)
  );
  bc_pe bc_pe_2 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_2_clock),
    .reset(bc_pe_2_reset),
    .io_ho_input(bc_pe_2_io_ho_input),
    .io_ve_input(bc_pe_2_io_ve_input),
    .io_input_valid(bc_pe_2_io_input_valid),
    .io_iormac(bc_pe_2_io_iormac),
    .io_ve_out(bc_pe_2_io_ve_out),
    .io_ho_out(bc_pe_2_io_ho_out),
    .io_res_out(bc_pe_2_io_res_out)
  );
  bc_pe bc_pe_3 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_3_clock),
    .reset(bc_pe_3_reset),
    .io_ho_input(bc_pe_3_io_ho_input),
    .io_ve_input(bc_pe_3_io_ve_input),
    .io_input_valid(bc_pe_3_io_input_valid),
    .io_iormac(bc_pe_3_io_iormac),
    .io_ve_out(bc_pe_3_io_ve_out),
    .io_ho_out(bc_pe_3_io_ho_out),
    .io_res_out(bc_pe_3_io_res_out)
  );
  bc_pe bc_pe_4 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_4_clock),
    .reset(bc_pe_4_reset),
    .io_ho_input(bc_pe_4_io_ho_input),
    .io_ve_input(bc_pe_4_io_ve_input),
    .io_input_valid(bc_pe_4_io_input_valid),
    .io_iormac(bc_pe_4_io_iormac),
    .io_ve_out(bc_pe_4_io_ve_out),
    .io_ho_out(bc_pe_4_io_ho_out),
    .io_res_out(bc_pe_4_io_res_out)
  );
  bc_pe bc_pe_5 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_5_clock),
    .reset(bc_pe_5_reset),
    .io_ho_input(bc_pe_5_io_ho_input),
    .io_ve_input(bc_pe_5_io_ve_input),
    .io_input_valid(bc_pe_5_io_input_valid),
    .io_iormac(bc_pe_5_io_iormac),
    .io_ve_out(bc_pe_5_io_ve_out),
    .io_ho_out(bc_pe_5_io_ho_out),
    .io_res_out(bc_pe_5_io_res_out)
  );
  bc_pe bc_pe_6 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_6_clock),
    .reset(bc_pe_6_reset),
    .io_ho_input(bc_pe_6_io_ho_input),
    .io_ve_input(bc_pe_6_io_ve_input),
    .io_input_valid(bc_pe_6_io_input_valid),
    .io_iormac(bc_pe_6_io_iormac),
    .io_ve_out(bc_pe_6_io_ve_out),
    .io_ho_out(bc_pe_6_io_ho_out),
    .io_res_out(bc_pe_6_io_res_out)
  );
  bc_pe bc_pe_7 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_7_clock),
    .reset(bc_pe_7_reset),
    .io_ho_input(bc_pe_7_io_ho_input),
    .io_ve_input(bc_pe_7_io_ve_input),
    .io_input_valid(bc_pe_7_io_input_valid),
    .io_iormac(bc_pe_7_io_iormac),
    .io_ve_out(bc_pe_7_io_ve_out),
    .io_ho_out(bc_pe_7_io_ho_out),
    .io_res_out(bc_pe_7_io_res_out)
  );
  bc_pe bc_pe_8 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_8_clock),
    .reset(bc_pe_8_reset),
    .io_ho_input(bc_pe_8_io_ho_input),
    .io_ve_input(bc_pe_8_io_ve_input),
    .io_input_valid(bc_pe_8_io_input_valid),
    .io_iormac(bc_pe_8_io_iormac),
    .io_ve_out(bc_pe_8_io_ve_out),
    .io_ho_out(bc_pe_8_io_ho_out),
    .io_res_out(bc_pe_8_io_res_out)
  );
  bc_pe bc_pe_9 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_9_clock),
    .reset(bc_pe_9_reset),
    .io_ho_input(bc_pe_9_io_ho_input),
    .io_ve_input(bc_pe_9_io_ve_input),
    .io_input_valid(bc_pe_9_io_input_valid),
    .io_iormac(bc_pe_9_io_iormac),
    .io_ve_out(bc_pe_9_io_ve_out),
    .io_ho_out(bc_pe_9_io_ho_out),
    .io_res_out(bc_pe_9_io_res_out)
  );
  bc_pe bc_pe_10 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_10_clock),
    .reset(bc_pe_10_reset),
    .io_ho_input(bc_pe_10_io_ho_input),
    .io_ve_input(bc_pe_10_io_ve_input),
    .io_input_valid(bc_pe_10_io_input_valid),
    .io_iormac(bc_pe_10_io_iormac),
    .io_ve_out(bc_pe_10_io_ve_out),
    .io_ho_out(bc_pe_10_io_ho_out),
    .io_res_out(bc_pe_10_io_res_out)
  );
  bc_pe bc_pe_11 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_11_clock),
    .reset(bc_pe_11_reset),
    .io_ho_input(bc_pe_11_io_ho_input),
    .io_ve_input(bc_pe_11_io_ve_input),
    .io_input_valid(bc_pe_11_io_input_valid),
    .io_iormac(bc_pe_11_io_iormac),
    .io_ve_out(bc_pe_11_io_ve_out),
    .io_ho_out(bc_pe_11_io_ho_out),
    .io_res_out(bc_pe_11_io_res_out)
  );
  bc_pe bc_pe_12 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_12_clock),
    .reset(bc_pe_12_reset),
    .io_ho_input(bc_pe_12_io_ho_input),
    .io_ve_input(bc_pe_12_io_ve_input),
    .io_input_valid(bc_pe_12_io_input_valid),
    .io_iormac(bc_pe_12_io_iormac),
    .io_ve_out(bc_pe_12_io_ve_out),
    .io_ho_out(bc_pe_12_io_ho_out),
    .io_res_out(bc_pe_12_io_res_out)
  );
  bc_pe bc_pe_13 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_13_clock),
    .reset(bc_pe_13_reset),
    .io_ho_input(bc_pe_13_io_ho_input),
    .io_ve_input(bc_pe_13_io_ve_input),
    .io_input_valid(bc_pe_13_io_input_valid),
    .io_iormac(bc_pe_13_io_iormac),
    .io_ve_out(bc_pe_13_io_ve_out),
    .io_ho_out(bc_pe_13_io_ho_out),
    .io_res_out(bc_pe_13_io_res_out)
  );
  bc_pe bc_pe_14 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_14_clock),
    .reset(bc_pe_14_reset),
    .io_ho_input(bc_pe_14_io_ho_input),
    .io_ve_input(bc_pe_14_io_ve_input),
    .io_input_valid(bc_pe_14_io_input_valid),
    .io_iormac(bc_pe_14_io_iormac),
    .io_ve_out(bc_pe_14_io_ve_out),
    .io_ho_out(bc_pe_14_io_ho_out),
    .io_res_out(bc_pe_14_io_res_out)
  );
  bc_pe bc_pe_15 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_15_clock),
    .reset(bc_pe_15_reset),
    .io_ho_input(bc_pe_15_io_ho_input),
    .io_ve_input(bc_pe_15_io_ve_input),
    .io_input_valid(bc_pe_15_io_input_valid),
    .io_iormac(bc_pe_15_io_iormac),
    .io_ve_out(bc_pe_15_io_ve_out),
    .io_ho_out(bc_pe_15_io_ho_out),
    .io_res_out(bc_pe_15_io_res_out)
  );
  bc_pe bc_pe_16 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_16_clock),
    .reset(bc_pe_16_reset),
    .io_ho_input(bc_pe_16_io_ho_input),
    .io_ve_input(bc_pe_16_io_ve_input),
    .io_input_valid(bc_pe_16_io_input_valid),
    .io_iormac(bc_pe_16_io_iormac),
    .io_ve_out(bc_pe_16_io_ve_out),
    .io_ho_out(bc_pe_16_io_ho_out),
    .io_res_out(bc_pe_16_io_res_out)
  );
  bc_pe bc_pe_17 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_17_clock),
    .reset(bc_pe_17_reset),
    .io_ho_input(bc_pe_17_io_ho_input),
    .io_ve_input(bc_pe_17_io_ve_input),
    .io_input_valid(bc_pe_17_io_input_valid),
    .io_iormac(bc_pe_17_io_iormac),
    .io_ve_out(bc_pe_17_io_ve_out),
    .io_ho_out(bc_pe_17_io_ho_out),
    .io_res_out(bc_pe_17_io_res_out)
  );
  bc_pe bc_pe_18 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_18_clock),
    .reset(bc_pe_18_reset),
    .io_ho_input(bc_pe_18_io_ho_input),
    .io_ve_input(bc_pe_18_io_ve_input),
    .io_input_valid(bc_pe_18_io_input_valid),
    .io_iormac(bc_pe_18_io_iormac),
    .io_ve_out(bc_pe_18_io_ve_out),
    .io_ho_out(bc_pe_18_io_ho_out),
    .io_res_out(bc_pe_18_io_res_out)
  );
  bc_pe bc_pe_19 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_19_clock),
    .reset(bc_pe_19_reset),
    .io_ho_input(bc_pe_19_io_ho_input),
    .io_ve_input(bc_pe_19_io_ve_input),
    .io_input_valid(bc_pe_19_io_input_valid),
    .io_iormac(bc_pe_19_io_iormac),
    .io_ve_out(bc_pe_19_io_ve_out),
    .io_ho_out(bc_pe_19_io_ho_out),
    .io_res_out(bc_pe_19_io_res_out)
  );
  bc_pe bc_pe_20 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_20_clock),
    .reset(bc_pe_20_reset),
    .io_ho_input(bc_pe_20_io_ho_input),
    .io_ve_input(bc_pe_20_io_ve_input),
    .io_input_valid(bc_pe_20_io_input_valid),
    .io_iormac(bc_pe_20_io_iormac),
    .io_ve_out(bc_pe_20_io_ve_out),
    .io_ho_out(bc_pe_20_io_ho_out),
    .io_res_out(bc_pe_20_io_res_out)
  );
  bc_pe bc_pe_21 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_21_clock),
    .reset(bc_pe_21_reset),
    .io_ho_input(bc_pe_21_io_ho_input),
    .io_ve_input(bc_pe_21_io_ve_input),
    .io_input_valid(bc_pe_21_io_input_valid),
    .io_iormac(bc_pe_21_io_iormac),
    .io_ve_out(bc_pe_21_io_ve_out),
    .io_ho_out(bc_pe_21_io_ho_out),
    .io_res_out(bc_pe_21_io_res_out)
  );
  bc_pe bc_pe_22 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_22_clock),
    .reset(bc_pe_22_reset),
    .io_ho_input(bc_pe_22_io_ho_input),
    .io_ve_input(bc_pe_22_io_ve_input),
    .io_input_valid(bc_pe_22_io_input_valid),
    .io_iormac(bc_pe_22_io_iormac),
    .io_ve_out(bc_pe_22_io_ve_out),
    .io_ho_out(bc_pe_22_io_ho_out),
    .io_res_out(bc_pe_22_io_res_out)
  );
  bc_pe bc_pe_23 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_23_clock),
    .reset(bc_pe_23_reset),
    .io_ho_input(bc_pe_23_io_ho_input),
    .io_ve_input(bc_pe_23_io_ve_input),
    .io_input_valid(bc_pe_23_io_input_valid),
    .io_iormac(bc_pe_23_io_iormac),
    .io_ve_out(bc_pe_23_io_ve_out),
    .io_ho_out(bc_pe_23_io_ho_out),
    .io_res_out(bc_pe_23_io_res_out)
  );
  bc_pe bc_pe_24 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_24_clock),
    .reset(bc_pe_24_reset),
    .io_ho_input(bc_pe_24_io_ho_input),
    .io_ve_input(bc_pe_24_io_ve_input),
    .io_input_valid(bc_pe_24_io_input_valid),
    .io_iormac(bc_pe_24_io_iormac),
    .io_ve_out(bc_pe_24_io_ve_out),
    .io_ho_out(bc_pe_24_io_ho_out),
    .io_res_out(bc_pe_24_io_res_out)
  );
  bc_pe bc_pe_25 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_25_clock),
    .reset(bc_pe_25_reset),
    .io_ho_input(bc_pe_25_io_ho_input),
    .io_ve_input(bc_pe_25_io_ve_input),
    .io_input_valid(bc_pe_25_io_input_valid),
    .io_iormac(bc_pe_25_io_iormac),
    .io_ve_out(bc_pe_25_io_ve_out),
    .io_ho_out(bc_pe_25_io_ho_out),
    .io_res_out(bc_pe_25_io_res_out)
  );
  bc_pe bc_pe_26 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_26_clock),
    .reset(bc_pe_26_reset),
    .io_ho_input(bc_pe_26_io_ho_input),
    .io_ve_input(bc_pe_26_io_ve_input),
    .io_input_valid(bc_pe_26_io_input_valid),
    .io_iormac(bc_pe_26_io_iormac),
    .io_ve_out(bc_pe_26_io_ve_out),
    .io_ho_out(bc_pe_26_io_ho_out),
    .io_res_out(bc_pe_26_io_res_out)
  );
  bc_pe bc_pe_27 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_27_clock),
    .reset(bc_pe_27_reset),
    .io_ho_input(bc_pe_27_io_ho_input),
    .io_ve_input(bc_pe_27_io_ve_input),
    .io_input_valid(bc_pe_27_io_input_valid),
    .io_iormac(bc_pe_27_io_iormac),
    .io_ve_out(bc_pe_27_io_ve_out),
    .io_ho_out(bc_pe_27_io_ho_out),
    .io_res_out(bc_pe_27_io_res_out)
  );
  bc_pe bc_pe_28 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_28_clock),
    .reset(bc_pe_28_reset),
    .io_ho_input(bc_pe_28_io_ho_input),
    .io_ve_input(bc_pe_28_io_ve_input),
    .io_input_valid(bc_pe_28_io_input_valid),
    .io_iormac(bc_pe_28_io_iormac),
    .io_ve_out(bc_pe_28_io_ve_out),
    .io_ho_out(bc_pe_28_io_ho_out),
    .io_res_out(bc_pe_28_io_res_out)
  );
  bc_pe bc_pe_29 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_29_clock),
    .reset(bc_pe_29_reset),
    .io_ho_input(bc_pe_29_io_ho_input),
    .io_ve_input(bc_pe_29_io_ve_input),
    .io_input_valid(bc_pe_29_io_input_valid),
    .io_iormac(bc_pe_29_io_iormac),
    .io_ve_out(bc_pe_29_io_ve_out),
    .io_ho_out(bc_pe_29_io_ho_out),
    .io_res_out(bc_pe_29_io_res_out)
  );
  bc_pe bc_pe_30 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_30_clock),
    .reset(bc_pe_30_reset),
    .io_ho_input(bc_pe_30_io_ho_input),
    .io_ve_input(bc_pe_30_io_ve_input),
    .io_input_valid(bc_pe_30_io_input_valid),
    .io_iormac(bc_pe_30_io_iormac),
    .io_ve_out(bc_pe_30_io_ve_out),
    .io_ho_out(bc_pe_30_io_ho_out),
    .io_res_out(bc_pe_30_io_res_out)
  );
  bc_pe bc_pe_31 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_31_clock),
    .reset(bc_pe_31_reset),
    .io_ho_input(bc_pe_31_io_ho_input),
    .io_ve_input(bc_pe_31_io_ve_input),
    .io_input_valid(bc_pe_31_io_input_valid),
    .io_iormac(bc_pe_31_io_iormac),
    .io_ve_out(bc_pe_31_io_ve_out),
    .io_ho_out(bc_pe_31_io_ho_out),
    .io_res_out(bc_pe_31_io_res_out)
  );
  bc_pe bc_pe_32 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_32_clock),
    .reset(bc_pe_32_reset),
    .io_ho_input(bc_pe_32_io_ho_input),
    .io_ve_input(bc_pe_32_io_ve_input),
    .io_input_valid(bc_pe_32_io_input_valid),
    .io_iormac(bc_pe_32_io_iormac),
    .io_ve_out(bc_pe_32_io_ve_out),
    .io_ho_out(bc_pe_32_io_ho_out),
    .io_res_out(bc_pe_32_io_res_out)
  );
  bc_pe bc_pe_33 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_33_clock),
    .reset(bc_pe_33_reset),
    .io_ho_input(bc_pe_33_io_ho_input),
    .io_ve_input(bc_pe_33_io_ve_input),
    .io_input_valid(bc_pe_33_io_input_valid),
    .io_iormac(bc_pe_33_io_iormac),
    .io_ve_out(bc_pe_33_io_ve_out),
    .io_ho_out(bc_pe_33_io_ho_out),
    .io_res_out(bc_pe_33_io_res_out)
  );
  bc_pe bc_pe_34 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_34_clock),
    .reset(bc_pe_34_reset),
    .io_ho_input(bc_pe_34_io_ho_input),
    .io_ve_input(bc_pe_34_io_ve_input),
    .io_input_valid(bc_pe_34_io_input_valid),
    .io_iormac(bc_pe_34_io_iormac),
    .io_ve_out(bc_pe_34_io_ve_out),
    .io_ho_out(bc_pe_34_io_ho_out),
    .io_res_out(bc_pe_34_io_res_out)
  );
  bc_pe bc_pe_35 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_35_clock),
    .reset(bc_pe_35_reset),
    .io_ho_input(bc_pe_35_io_ho_input),
    .io_ve_input(bc_pe_35_io_ve_input),
    .io_input_valid(bc_pe_35_io_input_valid),
    .io_iormac(bc_pe_35_io_iormac),
    .io_ve_out(bc_pe_35_io_ve_out),
    .io_ho_out(bc_pe_35_io_ho_out),
    .io_res_out(bc_pe_35_io_res_out)
  );
  bc_pe bc_pe_36 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_36_clock),
    .reset(bc_pe_36_reset),
    .io_ho_input(bc_pe_36_io_ho_input),
    .io_ve_input(bc_pe_36_io_ve_input),
    .io_input_valid(bc_pe_36_io_input_valid),
    .io_iormac(bc_pe_36_io_iormac),
    .io_ve_out(bc_pe_36_io_ve_out),
    .io_ho_out(bc_pe_36_io_ho_out),
    .io_res_out(bc_pe_36_io_res_out)
  );
  bc_pe bc_pe_37 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_37_clock),
    .reset(bc_pe_37_reset),
    .io_ho_input(bc_pe_37_io_ho_input),
    .io_ve_input(bc_pe_37_io_ve_input),
    .io_input_valid(bc_pe_37_io_input_valid),
    .io_iormac(bc_pe_37_io_iormac),
    .io_ve_out(bc_pe_37_io_ve_out),
    .io_ho_out(bc_pe_37_io_ho_out),
    .io_res_out(bc_pe_37_io_res_out)
  );
  bc_pe bc_pe_38 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_38_clock),
    .reset(bc_pe_38_reset),
    .io_ho_input(bc_pe_38_io_ho_input),
    .io_ve_input(bc_pe_38_io_ve_input),
    .io_input_valid(bc_pe_38_io_input_valid),
    .io_iormac(bc_pe_38_io_iormac),
    .io_ve_out(bc_pe_38_io_ve_out),
    .io_ho_out(bc_pe_38_io_ho_out),
    .io_res_out(bc_pe_38_io_res_out)
  );
  bc_pe bc_pe_39 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_39_clock),
    .reset(bc_pe_39_reset),
    .io_ho_input(bc_pe_39_io_ho_input),
    .io_ve_input(bc_pe_39_io_ve_input),
    .io_input_valid(bc_pe_39_io_input_valid),
    .io_iormac(bc_pe_39_io_iormac),
    .io_ve_out(bc_pe_39_io_ve_out),
    .io_ho_out(bc_pe_39_io_ho_out),
    .io_res_out(bc_pe_39_io_res_out)
  );
  bc_pe bc_pe_40 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_40_clock),
    .reset(bc_pe_40_reset),
    .io_ho_input(bc_pe_40_io_ho_input),
    .io_ve_input(bc_pe_40_io_ve_input),
    .io_input_valid(bc_pe_40_io_input_valid),
    .io_iormac(bc_pe_40_io_iormac),
    .io_ve_out(bc_pe_40_io_ve_out),
    .io_ho_out(bc_pe_40_io_ho_out),
    .io_res_out(bc_pe_40_io_res_out)
  );
  bc_pe bc_pe_41 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_41_clock),
    .reset(bc_pe_41_reset),
    .io_ho_input(bc_pe_41_io_ho_input),
    .io_ve_input(bc_pe_41_io_ve_input),
    .io_input_valid(bc_pe_41_io_input_valid),
    .io_iormac(bc_pe_41_io_iormac),
    .io_ve_out(bc_pe_41_io_ve_out),
    .io_ho_out(bc_pe_41_io_ho_out),
    .io_res_out(bc_pe_41_io_res_out)
  );
  bc_pe bc_pe_42 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_42_clock),
    .reset(bc_pe_42_reset),
    .io_ho_input(bc_pe_42_io_ho_input),
    .io_ve_input(bc_pe_42_io_ve_input),
    .io_input_valid(bc_pe_42_io_input_valid),
    .io_iormac(bc_pe_42_io_iormac),
    .io_ve_out(bc_pe_42_io_ve_out),
    .io_ho_out(bc_pe_42_io_ho_out),
    .io_res_out(bc_pe_42_io_res_out)
  );
  bc_pe bc_pe_43 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_43_clock),
    .reset(bc_pe_43_reset),
    .io_ho_input(bc_pe_43_io_ho_input),
    .io_ve_input(bc_pe_43_io_ve_input),
    .io_input_valid(bc_pe_43_io_input_valid),
    .io_iormac(bc_pe_43_io_iormac),
    .io_ve_out(bc_pe_43_io_ve_out),
    .io_ho_out(bc_pe_43_io_ho_out),
    .io_res_out(bc_pe_43_io_res_out)
  );
  bc_pe bc_pe_44 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_44_clock),
    .reset(bc_pe_44_reset),
    .io_ho_input(bc_pe_44_io_ho_input),
    .io_ve_input(bc_pe_44_io_ve_input),
    .io_input_valid(bc_pe_44_io_input_valid),
    .io_iormac(bc_pe_44_io_iormac),
    .io_ve_out(bc_pe_44_io_ve_out),
    .io_ho_out(bc_pe_44_io_ho_out),
    .io_res_out(bc_pe_44_io_res_out)
  );
  bc_pe bc_pe_45 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_45_clock),
    .reset(bc_pe_45_reset),
    .io_ho_input(bc_pe_45_io_ho_input),
    .io_ve_input(bc_pe_45_io_ve_input),
    .io_input_valid(bc_pe_45_io_input_valid),
    .io_iormac(bc_pe_45_io_iormac),
    .io_ve_out(bc_pe_45_io_ve_out),
    .io_ho_out(bc_pe_45_io_ho_out),
    .io_res_out(bc_pe_45_io_res_out)
  );
  bc_pe bc_pe_46 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_46_clock),
    .reset(bc_pe_46_reset),
    .io_ho_input(bc_pe_46_io_ho_input),
    .io_ve_input(bc_pe_46_io_ve_input),
    .io_input_valid(bc_pe_46_io_input_valid),
    .io_iormac(bc_pe_46_io_iormac),
    .io_ve_out(bc_pe_46_io_ve_out),
    .io_ho_out(bc_pe_46_io_ho_out),
    .io_res_out(bc_pe_46_io_res_out)
  );
  bc_pe bc_pe_47 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_47_clock),
    .reset(bc_pe_47_reset),
    .io_ho_input(bc_pe_47_io_ho_input),
    .io_ve_input(bc_pe_47_io_ve_input),
    .io_input_valid(bc_pe_47_io_input_valid),
    .io_iormac(bc_pe_47_io_iormac),
    .io_ve_out(bc_pe_47_io_ve_out),
    .io_ho_out(bc_pe_47_io_ho_out),
    .io_res_out(bc_pe_47_io_res_out)
  );
  bc_pe bc_pe_48 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_48_clock),
    .reset(bc_pe_48_reset),
    .io_ho_input(bc_pe_48_io_ho_input),
    .io_ve_input(bc_pe_48_io_ve_input),
    .io_input_valid(bc_pe_48_io_input_valid),
    .io_iormac(bc_pe_48_io_iormac),
    .io_ve_out(bc_pe_48_io_ve_out),
    .io_ho_out(bc_pe_48_io_ho_out),
    .io_res_out(bc_pe_48_io_res_out)
  );
  bc_pe bc_pe_49 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_49_clock),
    .reset(bc_pe_49_reset),
    .io_ho_input(bc_pe_49_io_ho_input),
    .io_ve_input(bc_pe_49_io_ve_input),
    .io_input_valid(bc_pe_49_io_input_valid),
    .io_iormac(bc_pe_49_io_iormac),
    .io_ve_out(bc_pe_49_io_ve_out),
    .io_ho_out(bc_pe_49_io_ho_out),
    .io_res_out(bc_pe_49_io_res_out)
  );
  bc_pe bc_pe_50 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_50_clock),
    .reset(bc_pe_50_reset),
    .io_ho_input(bc_pe_50_io_ho_input),
    .io_ve_input(bc_pe_50_io_ve_input),
    .io_input_valid(bc_pe_50_io_input_valid),
    .io_iormac(bc_pe_50_io_iormac),
    .io_ve_out(bc_pe_50_io_ve_out),
    .io_ho_out(bc_pe_50_io_ho_out),
    .io_res_out(bc_pe_50_io_res_out)
  );
  bc_pe bc_pe_51 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_51_clock),
    .reset(bc_pe_51_reset),
    .io_ho_input(bc_pe_51_io_ho_input),
    .io_ve_input(bc_pe_51_io_ve_input),
    .io_input_valid(bc_pe_51_io_input_valid),
    .io_iormac(bc_pe_51_io_iormac),
    .io_ve_out(bc_pe_51_io_ve_out),
    .io_ho_out(bc_pe_51_io_ho_out),
    .io_res_out(bc_pe_51_io_res_out)
  );
  bc_pe bc_pe_52 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_52_clock),
    .reset(bc_pe_52_reset),
    .io_ho_input(bc_pe_52_io_ho_input),
    .io_ve_input(bc_pe_52_io_ve_input),
    .io_input_valid(bc_pe_52_io_input_valid),
    .io_iormac(bc_pe_52_io_iormac),
    .io_ve_out(bc_pe_52_io_ve_out),
    .io_ho_out(bc_pe_52_io_ho_out),
    .io_res_out(bc_pe_52_io_res_out)
  );
  bc_pe bc_pe_53 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_53_clock),
    .reset(bc_pe_53_reset),
    .io_ho_input(bc_pe_53_io_ho_input),
    .io_ve_input(bc_pe_53_io_ve_input),
    .io_input_valid(bc_pe_53_io_input_valid),
    .io_iormac(bc_pe_53_io_iormac),
    .io_ve_out(bc_pe_53_io_ve_out),
    .io_ho_out(bc_pe_53_io_ho_out),
    .io_res_out(bc_pe_53_io_res_out)
  );
  bc_pe bc_pe_54 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_54_clock),
    .reset(bc_pe_54_reset),
    .io_ho_input(bc_pe_54_io_ho_input),
    .io_ve_input(bc_pe_54_io_ve_input),
    .io_input_valid(bc_pe_54_io_input_valid),
    .io_iormac(bc_pe_54_io_iormac),
    .io_ve_out(bc_pe_54_io_ve_out),
    .io_ho_out(bc_pe_54_io_ho_out),
    .io_res_out(bc_pe_54_io_res_out)
  );
  bc_pe bc_pe_55 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_55_clock),
    .reset(bc_pe_55_reset),
    .io_ho_input(bc_pe_55_io_ho_input),
    .io_ve_input(bc_pe_55_io_ve_input),
    .io_input_valid(bc_pe_55_io_input_valid),
    .io_iormac(bc_pe_55_io_iormac),
    .io_ve_out(bc_pe_55_io_ve_out),
    .io_ho_out(bc_pe_55_io_ho_out),
    .io_res_out(bc_pe_55_io_res_out)
  );
  bc_pe bc_pe_56 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_56_clock),
    .reset(bc_pe_56_reset),
    .io_ho_input(bc_pe_56_io_ho_input),
    .io_ve_input(bc_pe_56_io_ve_input),
    .io_input_valid(bc_pe_56_io_input_valid),
    .io_iormac(bc_pe_56_io_iormac),
    .io_ve_out(bc_pe_56_io_ve_out),
    .io_ho_out(bc_pe_56_io_ho_out),
    .io_res_out(bc_pe_56_io_res_out)
  );
  bc_pe bc_pe_57 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_57_clock),
    .reset(bc_pe_57_reset),
    .io_ho_input(bc_pe_57_io_ho_input),
    .io_ve_input(bc_pe_57_io_ve_input),
    .io_input_valid(bc_pe_57_io_input_valid),
    .io_iormac(bc_pe_57_io_iormac),
    .io_ve_out(bc_pe_57_io_ve_out),
    .io_ho_out(bc_pe_57_io_ho_out),
    .io_res_out(bc_pe_57_io_res_out)
  );
  bc_pe bc_pe_58 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_58_clock),
    .reset(bc_pe_58_reset),
    .io_ho_input(bc_pe_58_io_ho_input),
    .io_ve_input(bc_pe_58_io_ve_input),
    .io_input_valid(bc_pe_58_io_input_valid),
    .io_iormac(bc_pe_58_io_iormac),
    .io_ve_out(bc_pe_58_io_ve_out),
    .io_ho_out(bc_pe_58_io_ho_out),
    .io_res_out(bc_pe_58_io_res_out)
  );
  bc_pe bc_pe_59 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_59_clock),
    .reset(bc_pe_59_reset),
    .io_ho_input(bc_pe_59_io_ho_input),
    .io_ve_input(bc_pe_59_io_ve_input),
    .io_input_valid(bc_pe_59_io_input_valid),
    .io_iormac(bc_pe_59_io_iormac),
    .io_ve_out(bc_pe_59_io_ve_out),
    .io_ho_out(bc_pe_59_io_ho_out),
    .io_res_out(bc_pe_59_io_res_out)
  );
  bc_pe bc_pe_60 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_60_clock),
    .reset(bc_pe_60_reset),
    .io_ho_input(bc_pe_60_io_ho_input),
    .io_ve_input(bc_pe_60_io_ve_input),
    .io_input_valid(bc_pe_60_io_input_valid),
    .io_iormac(bc_pe_60_io_iormac),
    .io_ve_out(bc_pe_60_io_ve_out),
    .io_ho_out(bc_pe_60_io_ho_out),
    .io_res_out(bc_pe_60_io_res_out)
  );
  bc_pe bc_pe_61 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_61_clock),
    .reset(bc_pe_61_reset),
    .io_ho_input(bc_pe_61_io_ho_input),
    .io_ve_input(bc_pe_61_io_ve_input),
    .io_input_valid(bc_pe_61_io_input_valid),
    .io_iormac(bc_pe_61_io_iormac),
    .io_ve_out(bc_pe_61_io_ve_out),
    .io_ho_out(bc_pe_61_io_ho_out),
    .io_res_out(bc_pe_61_io_res_out)
  );
  bc_pe bc_pe_62 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_62_clock),
    .reset(bc_pe_62_reset),
    .io_ho_input(bc_pe_62_io_ho_input),
    .io_ve_input(bc_pe_62_io_ve_input),
    .io_input_valid(bc_pe_62_io_input_valid),
    .io_iormac(bc_pe_62_io_iormac),
    .io_ve_out(bc_pe_62_io_ve_out),
    .io_ho_out(bc_pe_62_io_ho_out),
    .io_res_out(bc_pe_62_io_res_out)
  );
  bc_pe bc_pe_63 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_63_clock),
    .reset(bc_pe_63_reset),
    .io_ho_input(bc_pe_63_io_ho_input),
    .io_ve_input(bc_pe_63_io_ve_input),
    .io_input_valid(bc_pe_63_io_input_valid),
    .io_iormac(bc_pe_63_io_iormac),
    .io_ve_out(bc_pe_63_io_ve_out),
    .io_ho_out(bc_pe_63_io_ho_out),
    .io_res_out(bc_pe_63_io_res_out)
  );
  bc_pe bc_pe_64 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_64_clock),
    .reset(bc_pe_64_reset),
    .io_ho_input(bc_pe_64_io_ho_input),
    .io_ve_input(bc_pe_64_io_ve_input),
    .io_input_valid(bc_pe_64_io_input_valid),
    .io_iormac(bc_pe_64_io_iormac),
    .io_ve_out(bc_pe_64_io_ve_out),
    .io_ho_out(bc_pe_64_io_ho_out),
    .io_res_out(bc_pe_64_io_res_out)
  );
  bc_pe bc_pe_65 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_65_clock),
    .reset(bc_pe_65_reset),
    .io_ho_input(bc_pe_65_io_ho_input),
    .io_ve_input(bc_pe_65_io_ve_input),
    .io_input_valid(bc_pe_65_io_input_valid),
    .io_iormac(bc_pe_65_io_iormac),
    .io_ve_out(bc_pe_65_io_ve_out),
    .io_ho_out(bc_pe_65_io_ho_out),
    .io_res_out(bc_pe_65_io_res_out)
  );
  bc_pe bc_pe_66 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_66_clock),
    .reset(bc_pe_66_reset),
    .io_ho_input(bc_pe_66_io_ho_input),
    .io_ve_input(bc_pe_66_io_ve_input),
    .io_input_valid(bc_pe_66_io_input_valid),
    .io_iormac(bc_pe_66_io_iormac),
    .io_ve_out(bc_pe_66_io_ve_out),
    .io_ho_out(bc_pe_66_io_ho_out),
    .io_res_out(bc_pe_66_io_res_out)
  );
  bc_pe bc_pe_67 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_67_clock),
    .reset(bc_pe_67_reset),
    .io_ho_input(bc_pe_67_io_ho_input),
    .io_ve_input(bc_pe_67_io_ve_input),
    .io_input_valid(bc_pe_67_io_input_valid),
    .io_iormac(bc_pe_67_io_iormac),
    .io_ve_out(bc_pe_67_io_ve_out),
    .io_ho_out(bc_pe_67_io_ho_out),
    .io_res_out(bc_pe_67_io_res_out)
  );
  bc_pe bc_pe_68 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_68_clock),
    .reset(bc_pe_68_reset),
    .io_ho_input(bc_pe_68_io_ho_input),
    .io_ve_input(bc_pe_68_io_ve_input),
    .io_input_valid(bc_pe_68_io_input_valid),
    .io_iormac(bc_pe_68_io_iormac),
    .io_ve_out(bc_pe_68_io_ve_out),
    .io_ho_out(bc_pe_68_io_ho_out),
    .io_res_out(bc_pe_68_io_res_out)
  );
  bc_pe bc_pe_69 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_69_clock),
    .reset(bc_pe_69_reset),
    .io_ho_input(bc_pe_69_io_ho_input),
    .io_ve_input(bc_pe_69_io_ve_input),
    .io_input_valid(bc_pe_69_io_input_valid),
    .io_iormac(bc_pe_69_io_iormac),
    .io_ve_out(bc_pe_69_io_ve_out),
    .io_ho_out(bc_pe_69_io_ho_out),
    .io_res_out(bc_pe_69_io_res_out)
  );
  bc_pe bc_pe_70 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_70_clock),
    .reset(bc_pe_70_reset),
    .io_ho_input(bc_pe_70_io_ho_input),
    .io_ve_input(bc_pe_70_io_ve_input),
    .io_input_valid(bc_pe_70_io_input_valid),
    .io_iormac(bc_pe_70_io_iormac),
    .io_ve_out(bc_pe_70_io_ve_out),
    .io_ho_out(bc_pe_70_io_ho_out),
    .io_res_out(bc_pe_70_io_res_out)
  );
  bc_pe bc_pe_71 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_71_clock),
    .reset(bc_pe_71_reset),
    .io_ho_input(bc_pe_71_io_ho_input),
    .io_ve_input(bc_pe_71_io_ve_input),
    .io_input_valid(bc_pe_71_io_input_valid),
    .io_iormac(bc_pe_71_io_iormac),
    .io_ve_out(bc_pe_71_io_ve_out),
    .io_ho_out(bc_pe_71_io_ho_out),
    .io_res_out(bc_pe_71_io_res_out)
  );
  bc_pe bc_pe_72 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_72_clock),
    .reset(bc_pe_72_reset),
    .io_ho_input(bc_pe_72_io_ho_input),
    .io_ve_input(bc_pe_72_io_ve_input),
    .io_input_valid(bc_pe_72_io_input_valid),
    .io_iormac(bc_pe_72_io_iormac),
    .io_ve_out(bc_pe_72_io_ve_out),
    .io_ho_out(bc_pe_72_io_ho_out),
    .io_res_out(bc_pe_72_io_res_out)
  );
  bc_pe bc_pe_73 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_73_clock),
    .reset(bc_pe_73_reset),
    .io_ho_input(bc_pe_73_io_ho_input),
    .io_ve_input(bc_pe_73_io_ve_input),
    .io_input_valid(bc_pe_73_io_input_valid),
    .io_iormac(bc_pe_73_io_iormac),
    .io_ve_out(bc_pe_73_io_ve_out),
    .io_ho_out(bc_pe_73_io_ho_out),
    .io_res_out(bc_pe_73_io_res_out)
  );
  bc_pe bc_pe_74 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_74_clock),
    .reset(bc_pe_74_reset),
    .io_ho_input(bc_pe_74_io_ho_input),
    .io_ve_input(bc_pe_74_io_ve_input),
    .io_input_valid(bc_pe_74_io_input_valid),
    .io_iormac(bc_pe_74_io_iormac),
    .io_ve_out(bc_pe_74_io_ve_out),
    .io_ho_out(bc_pe_74_io_ho_out),
    .io_res_out(bc_pe_74_io_res_out)
  );
  bc_pe bc_pe_75 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_75_clock),
    .reset(bc_pe_75_reset),
    .io_ho_input(bc_pe_75_io_ho_input),
    .io_ve_input(bc_pe_75_io_ve_input),
    .io_input_valid(bc_pe_75_io_input_valid),
    .io_iormac(bc_pe_75_io_iormac),
    .io_ve_out(bc_pe_75_io_ve_out),
    .io_ho_out(bc_pe_75_io_ho_out),
    .io_res_out(bc_pe_75_io_res_out)
  );
  bc_pe bc_pe_76 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_76_clock),
    .reset(bc_pe_76_reset),
    .io_ho_input(bc_pe_76_io_ho_input),
    .io_ve_input(bc_pe_76_io_ve_input),
    .io_input_valid(bc_pe_76_io_input_valid),
    .io_iormac(bc_pe_76_io_iormac),
    .io_ve_out(bc_pe_76_io_ve_out),
    .io_ho_out(bc_pe_76_io_ho_out),
    .io_res_out(bc_pe_76_io_res_out)
  );
  bc_pe bc_pe_77 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_77_clock),
    .reset(bc_pe_77_reset),
    .io_ho_input(bc_pe_77_io_ho_input),
    .io_ve_input(bc_pe_77_io_ve_input),
    .io_input_valid(bc_pe_77_io_input_valid),
    .io_iormac(bc_pe_77_io_iormac),
    .io_ve_out(bc_pe_77_io_ve_out),
    .io_ho_out(bc_pe_77_io_ho_out),
    .io_res_out(bc_pe_77_io_res_out)
  );
  bc_pe bc_pe_78 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_78_clock),
    .reset(bc_pe_78_reset),
    .io_ho_input(bc_pe_78_io_ho_input),
    .io_ve_input(bc_pe_78_io_ve_input),
    .io_input_valid(bc_pe_78_io_input_valid),
    .io_iormac(bc_pe_78_io_iormac),
    .io_ve_out(bc_pe_78_io_ve_out),
    .io_ho_out(bc_pe_78_io_ho_out),
    .io_res_out(bc_pe_78_io_res_out)
  );
  bc_pe bc_pe_79 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_79_clock),
    .reset(bc_pe_79_reset),
    .io_ho_input(bc_pe_79_io_ho_input),
    .io_ve_input(bc_pe_79_io_ve_input),
    .io_input_valid(bc_pe_79_io_input_valid),
    .io_iormac(bc_pe_79_io_iormac),
    .io_ve_out(bc_pe_79_io_ve_out),
    .io_ho_out(bc_pe_79_io_ho_out),
    .io_res_out(bc_pe_79_io_res_out)
  );
  bc_pe bc_pe_80 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_80_clock),
    .reset(bc_pe_80_reset),
    .io_ho_input(bc_pe_80_io_ho_input),
    .io_ve_input(bc_pe_80_io_ve_input),
    .io_input_valid(bc_pe_80_io_input_valid),
    .io_iormac(bc_pe_80_io_iormac),
    .io_ve_out(bc_pe_80_io_ve_out),
    .io_ho_out(bc_pe_80_io_ho_out),
    .io_res_out(bc_pe_80_io_res_out)
  );
  bc_pe bc_pe_81 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_81_clock),
    .reset(bc_pe_81_reset),
    .io_ho_input(bc_pe_81_io_ho_input),
    .io_ve_input(bc_pe_81_io_ve_input),
    .io_input_valid(bc_pe_81_io_input_valid),
    .io_iormac(bc_pe_81_io_iormac),
    .io_ve_out(bc_pe_81_io_ve_out),
    .io_ho_out(bc_pe_81_io_ho_out),
    .io_res_out(bc_pe_81_io_res_out)
  );
  bc_pe bc_pe_82 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_82_clock),
    .reset(bc_pe_82_reset),
    .io_ho_input(bc_pe_82_io_ho_input),
    .io_ve_input(bc_pe_82_io_ve_input),
    .io_input_valid(bc_pe_82_io_input_valid),
    .io_iormac(bc_pe_82_io_iormac),
    .io_ve_out(bc_pe_82_io_ve_out),
    .io_ho_out(bc_pe_82_io_ho_out),
    .io_res_out(bc_pe_82_io_res_out)
  );
  bc_pe bc_pe_83 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_83_clock),
    .reset(bc_pe_83_reset),
    .io_ho_input(bc_pe_83_io_ho_input),
    .io_ve_input(bc_pe_83_io_ve_input),
    .io_input_valid(bc_pe_83_io_input_valid),
    .io_iormac(bc_pe_83_io_iormac),
    .io_ve_out(bc_pe_83_io_ve_out),
    .io_ho_out(bc_pe_83_io_ho_out),
    .io_res_out(bc_pe_83_io_res_out)
  );
  bc_pe bc_pe_84 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_84_clock),
    .reset(bc_pe_84_reset),
    .io_ho_input(bc_pe_84_io_ho_input),
    .io_ve_input(bc_pe_84_io_ve_input),
    .io_input_valid(bc_pe_84_io_input_valid),
    .io_iormac(bc_pe_84_io_iormac),
    .io_ve_out(bc_pe_84_io_ve_out),
    .io_ho_out(bc_pe_84_io_ho_out),
    .io_res_out(bc_pe_84_io_res_out)
  );
  bc_pe bc_pe_85 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_85_clock),
    .reset(bc_pe_85_reset),
    .io_ho_input(bc_pe_85_io_ho_input),
    .io_ve_input(bc_pe_85_io_ve_input),
    .io_input_valid(bc_pe_85_io_input_valid),
    .io_iormac(bc_pe_85_io_iormac),
    .io_ve_out(bc_pe_85_io_ve_out),
    .io_ho_out(bc_pe_85_io_ho_out),
    .io_res_out(bc_pe_85_io_res_out)
  );
  bc_pe bc_pe_86 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_86_clock),
    .reset(bc_pe_86_reset),
    .io_ho_input(bc_pe_86_io_ho_input),
    .io_ve_input(bc_pe_86_io_ve_input),
    .io_input_valid(bc_pe_86_io_input_valid),
    .io_iormac(bc_pe_86_io_iormac),
    .io_ve_out(bc_pe_86_io_ve_out),
    .io_ho_out(bc_pe_86_io_ho_out),
    .io_res_out(bc_pe_86_io_res_out)
  );
  bc_pe bc_pe_87 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_87_clock),
    .reset(bc_pe_87_reset),
    .io_ho_input(bc_pe_87_io_ho_input),
    .io_ve_input(bc_pe_87_io_ve_input),
    .io_input_valid(bc_pe_87_io_input_valid),
    .io_iormac(bc_pe_87_io_iormac),
    .io_ve_out(bc_pe_87_io_ve_out),
    .io_ho_out(bc_pe_87_io_ho_out),
    .io_res_out(bc_pe_87_io_res_out)
  );
  bc_pe bc_pe_88 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_88_clock),
    .reset(bc_pe_88_reset),
    .io_ho_input(bc_pe_88_io_ho_input),
    .io_ve_input(bc_pe_88_io_ve_input),
    .io_input_valid(bc_pe_88_io_input_valid),
    .io_iormac(bc_pe_88_io_iormac),
    .io_ve_out(bc_pe_88_io_ve_out),
    .io_ho_out(bc_pe_88_io_ho_out),
    .io_res_out(bc_pe_88_io_res_out)
  );
  bc_pe bc_pe_89 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_89_clock),
    .reset(bc_pe_89_reset),
    .io_ho_input(bc_pe_89_io_ho_input),
    .io_ve_input(bc_pe_89_io_ve_input),
    .io_input_valid(bc_pe_89_io_input_valid),
    .io_iormac(bc_pe_89_io_iormac),
    .io_ve_out(bc_pe_89_io_ve_out),
    .io_ho_out(bc_pe_89_io_ho_out),
    .io_res_out(bc_pe_89_io_res_out)
  );
  bc_pe bc_pe_90 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_90_clock),
    .reset(bc_pe_90_reset),
    .io_ho_input(bc_pe_90_io_ho_input),
    .io_ve_input(bc_pe_90_io_ve_input),
    .io_input_valid(bc_pe_90_io_input_valid),
    .io_iormac(bc_pe_90_io_iormac),
    .io_ve_out(bc_pe_90_io_ve_out),
    .io_ho_out(bc_pe_90_io_ho_out),
    .io_res_out(bc_pe_90_io_res_out)
  );
  bc_pe bc_pe_91 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_91_clock),
    .reset(bc_pe_91_reset),
    .io_ho_input(bc_pe_91_io_ho_input),
    .io_ve_input(bc_pe_91_io_ve_input),
    .io_input_valid(bc_pe_91_io_input_valid),
    .io_iormac(bc_pe_91_io_iormac),
    .io_ve_out(bc_pe_91_io_ve_out),
    .io_ho_out(bc_pe_91_io_ho_out),
    .io_res_out(bc_pe_91_io_res_out)
  );
  bc_pe bc_pe_92 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_92_clock),
    .reset(bc_pe_92_reset),
    .io_ho_input(bc_pe_92_io_ho_input),
    .io_ve_input(bc_pe_92_io_ve_input),
    .io_input_valid(bc_pe_92_io_input_valid),
    .io_iormac(bc_pe_92_io_iormac),
    .io_ve_out(bc_pe_92_io_ve_out),
    .io_ho_out(bc_pe_92_io_ho_out),
    .io_res_out(bc_pe_92_io_res_out)
  );
  bc_pe bc_pe_93 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_93_clock),
    .reset(bc_pe_93_reset),
    .io_ho_input(bc_pe_93_io_ho_input),
    .io_ve_input(bc_pe_93_io_ve_input),
    .io_input_valid(bc_pe_93_io_input_valid),
    .io_iormac(bc_pe_93_io_iormac),
    .io_ve_out(bc_pe_93_io_ve_out),
    .io_ho_out(bc_pe_93_io_ho_out),
    .io_res_out(bc_pe_93_io_res_out)
  );
  bc_pe bc_pe_94 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_94_clock),
    .reset(bc_pe_94_reset),
    .io_ho_input(bc_pe_94_io_ho_input),
    .io_ve_input(bc_pe_94_io_ve_input),
    .io_input_valid(bc_pe_94_io_input_valid),
    .io_iormac(bc_pe_94_io_iormac),
    .io_ve_out(bc_pe_94_io_ve_out),
    .io_ho_out(bc_pe_94_io_ho_out),
    .io_res_out(bc_pe_94_io_res_out)
  );
  bc_pe bc_pe_95 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_95_clock),
    .reset(bc_pe_95_reset),
    .io_ho_input(bc_pe_95_io_ho_input),
    .io_ve_input(bc_pe_95_io_ve_input),
    .io_input_valid(bc_pe_95_io_input_valid),
    .io_iormac(bc_pe_95_io_iormac),
    .io_ve_out(bc_pe_95_io_ve_out),
    .io_ho_out(bc_pe_95_io_ho_out),
    .io_res_out(bc_pe_95_io_res_out)
  );
  bc_pe bc_pe_96 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_96_clock),
    .reset(bc_pe_96_reset),
    .io_ho_input(bc_pe_96_io_ho_input),
    .io_ve_input(bc_pe_96_io_ve_input),
    .io_input_valid(bc_pe_96_io_input_valid),
    .io_iormac(bc_pe_96_io_iormac),
    .io_ve_out(bc_pe_96_io_ve_out),
    .io_ho_out(bc_pe_96_io_ho_out),
    .io_res_out(bc_pe_96_io_res_out)
  );
  bc_pe bc_pe_97 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_97_clock),
    .reset(bc_pe_97_reset),
    .io_ho_input(bc_pe_97_io_ho_input),
    .io_ve_input(bc_pe_97_io_ve_input),
    .io_input_valid(bc_pe_97_io_input_valid),
    .io_iormac(bc_pe_97_io_iormac),
    .io_ve_out(bc_pe_97_io_ve_out),
    .io_ho_out(bc_pe_97_io_ho_out),
    .io_res_out(bc_pe_97_io_res_out)
  );
  bc_pe bc_pe_98 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_98_clock),
    .reset(bc_pe_98_reset),
    .io_ho_input(bc_pe_98_io_ho_input),
    .io_ve_input(bc_pe_98_io_ve_input),
    .io_input_valid(bc_pe_98_io_input_valid),
    .io_iormac(bc_pe_98_io_iormac),
    .io_ve_out(bc_pe_98_io_ve_out),
    .io_ho_out(bc_pe_98_io_ho_out),
    .io_res_out(bc_pe_98_io_res_out)
  );
  bc_pe bc_pe_99 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_99_clock),
    .reset(bc_pe_99_reset),
    .io_ho_input(bc_pe_99_io_ho_input),
    .io_ve_input(bc_pe_99_io_ve_input),
    .io_input_valid(bc_pe_99_io_input_valid),
    .io_iormac(bc_pe_99_io_iormac),
    .io_ve_out(bc_pe_99_io_ve_out),
    .io_ho_out(bc_pe_99_io_ho_out),
    .io_res_out(bc_pe_99_io_res_out)
  );
  bc_pe bc_pe_100 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_100_clock),
    .reset(bc_pe_100_reset),
    .io_ho_input(bc_pe_100_io_ho_input),
    .io_ve_input(bc_pe_100_io_ve_input),
    .io_input_valid(bc_pe_100_io_input_valid),
    .io_iormac(bc_pe_100_io_iormac),
    .io_ve_out(bc_pe_100_io_ve_out),
    .io_ho_out(bc_pe_100_io_ho_out),
    .io_res_out(bc_pe_100_io_res_out)
  );
  bc_pe bc_pe_101 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_101_clock),
    .reset(bc_pe_101_reset),
    .io_ho_input(bc_pe_101_io_ho_input),
    .io_ve_input(bc_pe_101_io_ve_input),
    .io_input_valid(bc_pe_101_io_input_valid),
    .io_iormac(bc_pe_101_io_iormac),
    .io_ve_out(bc_pe_101_io_ve_out),
    .io_ho_out(bc_pe_101_io_ho_out),
    .io_res_out(bc_pe_101_io_res_out)
  );
  bc_pe bc_pe_102 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_102_clock),
    .reset(bc_pe_102_reset),
    .io_ho_input(bc_pe_102_io_ho_input),
    .io_ve_input(bc_pe_102_io_ve_input),
    .io_input_valid(bc_pe_102_io_input_valid),
    .io_iormac(bc_pe_102_io_iormac),
    .io_ve_out(bc_pe_102_io_ve_out),
    .io_ho_out(bc_pe_102_io_ho_out),
    .io_res_out(bc_pe_102_io_res_out)
  );
  bc_pe bc_pe_103 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_103_clock),
    .reset(bc_pe_103_reset),
    .io_ho_input(bc_pe_103_io_ho_input),
    .io_ve_input(bc_pe_103_io_ve_input),
    .io_input_valid(bc_pe_103_io_input_valid),
    .io_iormac(bc_pe_103_io_iormac),
    .io_ve_out(bc_pe_103_io_ve_out),
    .io_ho_out(bc_pe_103_io_ho_out),
    .io_res_out(bc_pe_103_io_res_out)
  );
  bc_pe bc_pe_104 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_104_clock),
    .reset(bc_pe_104_reset),
    .io_ho_input(bc_pe_104_io_ho_input),
    .io_ve_input(bc_pe_104_io_ve_input),
    .io_input_valid(bc_pe_104_io_input_valid),
    .io_iormac(bc_pe_104_io_iormac),
    .io_ve_out(bc_pe_104_io_ve_out),
    .io_ho_out(bc_pe_104_io_ho_out),
    .io_res_out(bc_pe_104_io_res_out)
  );
  bc_pe bc_pe_105 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_105_clock),
    .reset(bc_pe_105_reset),
    .io_ho_input(bc_pe_105_io_ho_input),
    .io_ve_input(bc_pe_105_io_ve_input),
    .io_input_valid(bc_pe_105_io_input_valid),
    .io_iormac(bc_pe_105_io_iormac),
    .io_ve_out(bc_pe_105_io_ve_out),
    .io_ho_out(bc_pe_105_io_ho_out),
    .io_res_out(bc_pe_105_io_res_out)
  );
  bc_pe bc_pe_106 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_106_clock),
    .reset(bc_pe_106_reset),
    .io_ho_input(bc_pe_106_io_ho_input),
    .io_ve_input(bc_pe_106_io_ve_input),
    .io_input_valid(bc_pe_106_io_input_valid),
    .io_iormac(bc_pe_106_io_iormac),
    .io_ve_out(bc_pe_106_io_ve_out),
    .io_ho_out(bc_pe_106_io_ho_out),
    .io_res_out(bc_pe_106_io_res_out)
  );
  bc_pe bc_pe_107 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_107_clock),
    .reset(bc_pe_107_reset),
    .io_ho_input(bc_pe_107_io_ho_input),
    .io_ve_input(bc_pe_107_io_ve_input),
    .io_input_valid(bc_pe_107_io_input_valid),
    .io_iormac(bc_pe_107_io_iormac),
    .io_ve_out(bc_pe_107_io_ve_out),
    .io_ho_out(bc_pe_107_io_ho_out),
    .io_res_out(bc_pe_107_io_res_out)
  );
  bc_pe bc_pe_108 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_108_clock),
    .reset(bc_pe_108_reset),
    .io_ho_input(bc_pe_108_io_ho_input),
    .io_ve_input(bc_pe_108_io_ve_input),
    .io_input_valid(bc_pe_108_io_input_valid),
    .io_iormac(bc_pe_108_io_iormac),
    .io_ve_out(bc_pe_108_io_ve_out),
    .io_ho_out(bc_pe_108_io_ho_out),
    .io_res_out(bc_pe_108_io_res_out)
  );
  bc_pe bc_pe_109 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_109_clock),
    .reset(bc_pe_109_reset),
    .io_ho_input(bc_pe_109_io_ho_input),
    .io_ve_input(bc_pe_109_io_ve_input),
    .io_input_valid(bc_pe_109_io_input_valid),
    .io_iormac(bc_pe_109_io_iormac),
    .io_ve_out(bc_pe_109_io_ve_out),
    .io_ho_out(bc_pe_109_io_ho_out),
    .io_res_out(bc_pe_109_io_res_out)
  );
  bc_pe bc_pe_110 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_110_clock),
    .reset(bc_pe_110_reset),
    .io_ho_input(bc_pe_110_io_ho_input),
    .io_ve_input(bc_pe_110_io_ve_input),
    .io_input_valid(bc_pe_110_io_input_valid),
    .io_iormac(bc_pe_110_io_iormac),
    .io_ve_out(bc_pe_110_io_ve_out),
    .io_ho_out(bc_pe_110_io_ho_out),
    .io_res_out(bc_pe_110_io_res_out)
  );
  bc_pe bc_pe_111 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_111_clock),
    .reset(bc_pe_111_reset),
    .io_ho_input(bc_pe_111_io_ho_input),
    .io_ve_input(bc_pe_111_io_ve_input),
    .io_input_valid(bc_pe_111_io_input_valid),
    .io_iormac(bc_pe_111_io_iormac),
    .io_ve_out(bc_pe_111_io_ve_out),
    .io_ho_out(bc_pe_111_io_ho_out),
    .io_res_out(bc_pe_111_io_res_out)
  );
  bc_pe bc_pe_112 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_112_clock),
    .reset(bc_pe_112_reset),
    .io_ho_input(bc_pe_112_io_ho_input),
    .io_ve_input(bc_pe_112_io_ve_input),
    .io_input_valid(bc_pe_112_io_input_valid),
    .io_iormac(bc_pe_112_io_iormac),
    .io_ve_out(bc_pe_112_io_ve_out),
    .io_ho_out(bc_pe_112_io_ho_out),
    .io_res_out(bc_pe_112_io_res_out)
  );
  bc_pe bc_pe_113 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_113_clock),
    .reset(bc_pe_113_reset),
    .io_ho_input(bc_pe_113_io_ho_input),
    .io_ve_input(bc_pe_113_io_ve_input),
    .io_input_valid(bc_pe_113_io_input_valid),
    .io_iormac(bc_pe_113_io_iormac),
    .io_ve_out(bc_pe_113_io_ve_out),
    .io_ho_out(bc_pe_113_io_ho_out),
    .io_res_out(bc_pe_113_io_res_out)
  );
  bc_pe bc_pe_114 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_114_clock),
    .reset(bc_pe_114_reset),
    .io_ho_input(bc_pe_114_io_ho_input),
    .io_ve_input(bc_pe_114_io_ve_input),
    .io_input_valid(bc_pe_114_io_input_valid),
    .io_iormac(bc_pe_114_io_iormac),
    .io_ve_out(bc_pe_114_io_ve_out),
    .io_ho_out(bc_pe_114_io_ho_out),
    .io_res_out(bc_pe_114_io_res_out)
  );
  bc_pe bc_pe_115 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_115_clock),
    .reset(bc_pe_115_reset),
    .io_ho_input(bc_pe_115_io_ho_input),
    .io_ve_input(bc_pe_115_io_ve_input),
    .io_input_valid(bc_pe_115_io_input_valid),
    .io_iormac(bc_pe_115_io_iormac),
    .io_ve_out(bc_pe_115_io_ve_out),
    .io_ho_out(bc_pe_115_io_ho_out),
    .io_res_out(bc_pe_115_io_res_out)
  );
  bc_pe bc_pe_116 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_116_clock),
    .reset(bc_pe_116_reset),
    .io_ho_input(bc_pe_116_io_ho_input),
    .io_ve_input(bc_pe_116_io_ve_input),
    .io_input_valid(bc_pe_116_io_input_valid),
    .io_iormac(bc_pe_116_io_iormac),
    .io_ve_out(bc_pe_116_io_ve_out),
    .io_ho_out(bc_pe_116_io_ho_out),
    .io_res_out(bc_pe_116_io_res_out)
  );
  bc_pe bc_pe_117 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_117_clock),
    .reset(bc_pe_117_reset),
    .io_ho_input(bc_pe_117_io_ho_input),
    .io_ve_input(bc_pe_117_io_ve_input),
    .io_input_valid(bc_pe_117_io_input_valid),
    .io_iormac(bc_pe_117_io_iormac),
    .io_ve_out(bc_pe_117_io_ve_out),
    .io_ho_out(bc_pe_117_io_ho_out),
    .io_res_out(bc_pe_117_io_res_out)
  );
  bc_pe bc_pe_118 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_118_clock),
    .reset(bc_pe_118_reset),
    .io_ho_input(bc_pe_118_io_ho_input),
    .io_ve_input(bc_pe_118_io_ve_input),
    .io_input_valid(bc_pe_118_io_input_valid),
    .io_iormac(bc_pe_118_io_iormac),
    .io_ve_out(bc_pe_118_io_ve_out),
    .io_ho_out(bc_pe_118_io_ho_out),
    .io_res_out(bc_pe_118_io_res_out)
  );
  bc_pe bc_pe_119 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_119_clock),
    .reset(bc_pe_119_reset),
    .io_ho_input(bc_pe_119_io_ho_input),
    .io_ve_input(bc_pe_119_io_ve_input),
    .io_input_valid(bc_pe_119_io_input_valid),
    .io_iormac(bc_pe_119_io_iormac),
    .io_ve_out(bc_pe_119_io_ve_out),
    .io_ho_out(bc_pe_119_io_ho_out),
    .io_res_out(bc_pe_119_io_res_out)
  );
  bc_pe bc_pe_120 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_120_clock),
    .reset(bc_pe_120_reset),
    .io_ho_input(bc_pe_120_io_ho_input),
    .io_ve_input(bc_pe_120_io_ve_input),
    .io_input_valid(bc_pe_120_io_input_valid),
    .io_iormac(bc_pe_120_io_iormac),
    .io_ve_out(bc_pe_120_io_ve_out),
    .io_ho_out(bc_pe_120_io_ho_out),
    .io_res_out(bc_pe_120_io_res_out)
  );
  bc_pe bc_pe_121 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_121_clock),
    .reset(bc_pe_121_reset),
    .io_ho_input(bc_pe_121_io_ho_input),
    .io_ve_input(bc_pe_121_io_ve_input),
    .io_input_valid(bc_pe_121_io_input_valid),
    .io_iormac(bc_pe_121_io_iormac),
    .io_ve_out(bc_pe_121_io_ve_out),
    .io_ho_out(bc_pe_121_io_ho_out),
    .io_res_out(bc_pe_121_io_res_out)
  );
  bc_pe bc_pe_122 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_122_clock),
    .reset(bc_pe_122_reset),
    .io_ho_input(bc_pe_122_io_ho_input),
    .io_ve_input(bc_pe_122_io_ve_input),
    .io_input_valid(bc_pe_122_io_input_valid),
    .io_iormac(bc_pe_122_io_iormac),
    .io_ve_out(bc_pe_122_io_ve_out),
    .io_ho_out(bc_pe_122_io_ho_out),
    .io_res_out(bc_pe_122_io_res_out)
  );
  bc_pe bc_pe_123 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_123_clock),
    .reset(bc_pe_123_reset),
    .io_ho_input(bc_pe_123_io_ho_input),
    .io_ve_input(bc_pe_123_io_ve_input),
    .io_input_valid(bc_pe_123_io_input_valid),
    .io_iormac(bc_pe_123_io_iormac),
    .io_ve_out(bc_pe_123_io_ve_out),
    .io_ho_out(bc_pe_123_io_ho_out),
    .io_res_out(bc_pe_123_io_res_out)
  );
  bc_pe bc_pe_124 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_124_clock),
    .reset(bc_pe_124_reset),
    .io_ho_input(bc_pe_124_io_ho_input),
    .io_ve_input(bc_pe_124_io_ve_input),
    .io_input_valid(bc_pe_124_io_input_valid),
    .io_iormac(bc_pe_124_io_iormac),
    .io_ve_out(bc_pe_124_io_ve_out),
    .io_ho_out(bc_pe_124_io_ho_out),
    .io_res_out(bc_pe_124_io_res_out)
  );
  bc_pe bc_pe_125 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_125_clock),
    .reset(bc_pe_125_reset),
    .io_ho_input(bc_pe_125_io_ho_input),
    .io_ve_input(bc_pe_125_io_ve_input),
    .io_input_valid(bc_pe_125_io_input_valid),
    .io_iormac(bc_pe_125_io_iormac),
    .io_ve_out(bc_pe_125_io_ve_out),
    .io_ho_out(bc_pe_125_io_ho_out),
    .io_res_out(bc_pe_125_io_res_out)
  );
  bc_pe bc_pe_126 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_126_clock),
    .reset(bc_pe_126_reset),
    .io_ho_input(bc_pe_126_io_ho_input),
    .io_ve_input(bc_pe_126_io_ve_input),
    .io_input_valid(bc_pe_126_io_input_valid),
    .io_iormac(bc_pe_126_io_iormac),
    .io_ve_out(bc_pe_126_io_ve_out),
    .io_ho_out(bc_pe_126_io_ho_out),
    .io_res_out(bc_pe_126_io_res_out)
  );
  bc_pe bc_pe_127 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_127_clock),
    .reset(bc_pe_127_reset),
    .io_ho_input(bc_pe_127_io_ho_input),
    .io_ve_input(bc_pe_127_io_ve_input),
    .io_input_valid(bc_pe_127_io_input_valid),
    .io_iormac(bc_pe_127_io_iormac),
    .io_ve_out(bc_pe_127_io_ve_out),
    .io_ho_out(bc_pe_127_io_ho_out),
    .io_res_out(bc_pe_127_io_res_out)
  );
  bc_pe bc_pe_128 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_128_clock),
    .reset(bc_pe_128_reset),
    .io_ho_input(bc_pe_128_io_ho_input),
    .io_ve_input(bc_pe_128_io_ve_input),
    .io_input_valid(bc_pe_128_io_input_valid),
    .io_iormac(bc_pe_128_io_iormac),
    .io_ve_out(bc_pe_128_io_ve_out),
    .io_ho_out(bc_pe_128_io_ho_out),
    .io_res_out(bc_pe_128_io_res_out)
  );
  bc_pe bc_pe_129 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_129_clock),
    .reset(bc_pe_129_reset),
    .io_ho_input(bc_pe_129_io_ho_input),
    .io_ve_input(bc_pe_129_io_ve_input),
    .io_input_valid(bc_pe_129_io_input_valid),
    .io_iormac(bc_pe_129_io_iormac),
    .io_ve_out(bc_pe_129_io_ve_out),
    .io_ho_out(bc_pe_129_io_ho_out),
    .io_res_out(bc_pe_129_io_res_out)
  );
  bc_pe bc_pe_130 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_130_clock),
    .reset(bc_pe_130_reset),
    .io_ho_input(bc_pe_130_io_ho_input),
    .io_ve_input(bc_pe_130_io_ve_input),
    .io_input_valid(bc_pe_130_io_input_valid),
    .io_iormac(bc_pe_130_io_iormac),
    .io_ve_out(bc_pe_130_io_ve_out),
    .io_ho_out(bc_pe_130_io_ho_out),
    .io_res_out(bc_pe_130_io_res_out)
  );
  bc_pe bc_pe_131 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_131_clock),
    .reset(bc_pe_131_reset),
    .io_ho_input(bc_pe_131_io_ho_input),
    .io_ve_input(bc_pe_131_io_ve_input),
    .io_input_valid(bc_pe_131_io_input_valid),
    .io_iormac(bc_pe_131_io_iormac),
    .io_ve_out(bc_pe_131_io_ve_out),
    .io_ho_out(bc_pe_131_io_ho_out),
    .io_res_out(bc_pe_131_io_res_out)
  );
  bc_pe bc_pe_132 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_132_clock),
    .reset(bc_pe_132_reset),
    .io_ho_input(bc_pe_132_io_ho_input),
    .io_ve_input(bc_pe_132_io_ve_input),
    .io_input_valid(bc_pe_132_io_input_valid),
    .io_iormac(bc_pe_132_io_iormac),
    .io_ve_out(bc_pe_132_io_ve_out),
    .io_ho_out(bc_pe_132_io_ho_out),
    .io_res_out(bc_pe_132_io_res_out)
  );
  bc_pe bc_pe_133 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_133_clock),
    .reset(bc_pe_133_reset),
    .io_ho_input(bc_pe_133_io_ho_input),
    .io_ve_input(bc_pe_133_io_ve_input),
    .io_input_valid(bc_pe_133_io_input_valid),
    .io_iormac(bc_pe_133_io_iormac),
    .io_ve_out(bc_pe_133_io_ve_out),
    .io_ho_out(bc_pe_133_io_ho_out),
    .io_res_out(bc_pe_133_io_res_out)
  );
  bc_pe bc_pe_134 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_134_clock),
    .reset(bc_pe_134_reset),
    .io_ho_input(bc_pe_134_io_ho_input),
    .io_ve_input(bc_pe_134_io_ve_input),
    .io_input_valid(bc_pe_134_io_input_valid),
    .io_iormac(bc_pe_134_io_iormac),
    .io_ve_out(bc_pe_134_io_ve_out),
    .io_ho_out(bc_pe_134_io_ho_out),
    .io_res_out(bc_pe_134_io_res_out)
  );
  bc_pe bc_pe_135 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_135_clock),
    .reset(bc_pe_135_reset),
    .io_ho_input(bc_pe_135_io_ho_input),
    .io_ve_input(bc_pe_135_io_ve_input),
    .io_input_valid(bc_pe_135_io_input_valid),
    .io_iormac(bc_pe_135_io_iormac),
    .io_ve_out(bc_pe_135_io_ve_out),
    .io_ho_out(bc_pe_135_io_ho_out),
    .io_res_out(bc_pe_135_io_res_out)
  );
  bc_pe bc_pe_136 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_136_clock),
    .reset(bc_pe_136_reset),
    .io_ho_input(bc_pe_136_io_ho_input),
    .io_ve_input(bc_pe_136_io_ve_input),
    .io_input_valid(bc_pe_136_io_input_valid),
    .io_iormac(bc_pe_136_io_iormac),
    .io_ve_out(bc_pe_136_io_ve_out),
    .io_ho_out(bc_pe_136_io_ho_out),
    .io_res_out(bc_pe_136_io_res_out)
  );
  bc_pe bc_pe_137 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_137_clock),
    .reset(bc_pe_137_reset),
    .io_ho_input(bc_pe_137_io_ho_input),
    .io_ve_input(bc_pe_137_io_ve_input),
    .io_input_valid(bc_pe_137_io_input_valid),
    .io_iormac(bc_pe_137_io_iormac),
    .io_ve_out(bc_pe_137_io_ve_out),
    .io_ho_out(bc_pe_137_io_ho_out),
    .io_res_out(bc_pe_137_io_res_out)
  );
  bc_pe bc_pe_138 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_138_clock),
    .reset(bc_pe_138_reset),
    .io_ho_input(bc_pe_138_io_ho_input),
    .io_ve_input(bc_pe_138_io_ve_input),
    .io_input_valid(bc_pe_138_io_input_valid),
    .io_iormac(bc_pe_138_io_iormac),
    .io_ve_out(bc_pe_138_io_ve_out),
    .io_ho_out(bc_pe_138_io_ho_out),
    .io_res_out(bc_pe_138_io_res_out)
  );
  bc_pe bc_pe_139 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_139_clock),
    .reset(bc_pe_139_reset),
    .io_ho_input(bc_pe_139_io_ho_input),
    .io_ve_input(bc_pe_139_io_ve_input),
    .io_input_valid(bc_pe_139_io_input_valid),
    .io_iormac(bc_pe_139_io_iormac),
    .io_ve_out(bc_pe_139_io_ve_out),
    .io_ho_out(bc_pe_139_io_ho_out),
    .io_res_out(bc_pe_139_io_res_out)
  );
  bc_pe bc_pe_140 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_140_clock),
    .reset(bc_pe_140_reset),
    .io_ho_input(bc_pe_140_io_ho_input),
    .io_ve_input(bc_pe_140_io_ve_input),
    .io_input_valid(bc_pe_140_io_input_valid),
    .io_iormac(bc_pe_140_io_iormac),
    .io_ve_out(bc_pe_140_io_ve_out),
    .io_ho_out(bc_pe_140_io_ho_out),
    .io_res_out(bc_pe_140_io_res_out)
  );
  bc_pe bc_pe_141 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_141_clock),
    .reset(bc_pe_141_reset),
    .io_ho_input(bc_pe_141_io_ho_input),
    .io_ve_input(bc_pe_141_io_ve_input),
    .io_input_valid(bc_pe_141_io_input_valid),
    .io_iormac(bc_pe_141_io_iormac),
    .io_ve_out(bc_pe_141_io_ve_out),
    .io_ho_out(bc_pe_141_io_ho_out),
    .io_res_out(bc_pe_141_io_res_out)
  );
  bc_pe bc_pe_142 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_142_clock),
    .reset(bc_pe_142_reset),
    .io_ho_input(bc_pe_142_io_ho_input),
    .io_ve_input(bc_pe_142_io_ve_input),
    .io_input_valid(bc_pe_142_io_input_valid),
    .io_iormac(bc_pe_142_io_iormac),
    .io_ve_out(bc_pe_142_io_ve_out),
    .io_ho_out(bc_pe_142_io_ho_out),
    .io_res_out(bc_pe_142_io_res_out)
  );
  bc_pe bc_pe_143 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_143_clock),
    .reset(bc_pe_143_reset),
    .io_ho_input(bc_pe_143_io_ho_input),
    .io_ve_input(bc_pe_143_io_ve_input),
    .io_input_valid(bc_pe_143_io_input_valid),
    .io_iormac(bc_pe_143_io_iormac),
    .io_ve_out(bc_pe_143_io_ve_out),
    .io_ho_out(bc_pe_143_io_ho_out),
    .io_res_out(bc_pe_143_io_res_out)
  );
  bc_pe bc_pe_144 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_144_clock),
    .reset(bc_pe_144_reset),
    .io_ho_input(bc_pe_144_io_ho_input),
    .io_ve_input(bc_pe_144_io_ve_input),
    .io_input_valid(bc_pe_144_io_input_valid),
    .io_iormac(bc_pe_144_io_iormac),
    .io_ve_out(bc_pe_144_io_ve_out),
    .io_ho_out(bc_pe_144_io_ho_out),
    .io_res_out(bc_pe_144_io_res_out)
  );
  bc_pe bc_pe_145 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_145_clock),
    .reset(bc_pe_145_reset),
    .io_ho_input(bc_pe_145_io_ho_input),
    .io_ve_input(bc_pe_145_io_ve_input),
    .io_input_valid(bc_pe_145_io_input_valid),
    .io_iormac(bc_pe_145_io_iormac),
    .io_ve_out(bc_pe_145_io_ve_out),
    .io_ho_out(bc_pe_145_io_ho_out),
    .io_res_out(bc_pe_145_io_res_out)
  );
  bc_pe bc_pe_146 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_146_clock),
    .reset(bc_pe_146_reset),
    .io_ho_input(bc_pe_146_io_ho_input),
    .io_ve_input(bc_pe_146_io_ve_input),
    .io_input_valid(bc_pe_146_io_input_valid),
    .io_iormac(bc_pe_146_io_iormac),
    .io_ve_out(bc_pe_146_io_ve_out),
    .io_ho_out(bc_pe_146_io_ho_out),
    .io_res_out(bc_pe_146_io_res_out)
  );
  bc_pe bc_pe_147 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_147_clock),
    .reset(bc_pe_147_reset),
    .io_ho_input(bc_pe_147_io_ho_input),
    .io_ve_input(bc_pe_147_io_ve_input),
    .io_input_valid(bc_pe_147_io_input_valid),
    .io_iormac(bc_pe_147_io_iormac),
    .io_ve_out(bc_pe_147_io_ve_out),
    .io_ho_out(bc_pe_147_io_ho_out),
    .io_res_out(bc_pe_147_io_res_out)
  );
  bc_pe bc_pe_148 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_148_clock),
    .reset(bc_pe_148_reset),
    .io_ho_input(bc_pe_148_io_ho_input),
    .io_ve_input(bc_pe_148_io_ve_input),
    .io_input_valid(bc_pe_148_io_input_valid),
    .io_iormac(bc_pe_148_io_iormac),
    .io_ve_out(bc_pe_148_io_ve_out),
    .io_ho_out(bc_pe_148_io_ho_out),
    .io_res_out(bc_pe_148_io_res_out)
  );
  bc_pe bc_pe_149 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_149_clock),
    .reset(bc_pe_149_reset),
    .io_ho_input(bc_pe_149_io_ho_input),
    .io_ve_input(bc_pe_149_io_ve_input),
    .io_input_valid(bc_pe_149_io_input_valid),
    .io_iormac(bc_pe_149_io_iormac),
    .io_ve_out(bc_pe_149_io_ve_out),
    .io_ho_out(bc_pe_149_io_ho_out),
    .io_res_out(bc_pe_149_io_res_out)
  );
  bc_pe bc_pe_150 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_150_clock),
    .reset(bc_pe_150_reset),
    .io_ho_input(bc_pe_150_io_ho_input),
    .io_ve_input(bc_pe_150_io_ve_input),
    .io_input_valid(bc_pe_150_io_input_valid),
    .io_iormac(bc_pe_150_io_iormac),
    .io_ve_out(bc_pe_150_io_ve_out),
    .io_ho_out(bc_pe_150_io_ho_out),
    .io_res_out(bc_pe_150_io_res_out)
  );
  bc_pe bc_pe_151 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_151_clock),
    .reset(bc_pe_151_reset),
    .io_ho_input(bc_pe_151_io_ho_input),
    .io_ve_input(bc_pe_151_io_ve_input),
    .io_input_valid(bc_pe_151_io_input_valid),
    .io_iormac(bc_pe_151_io_iormac),
    .io_ve_out(bc_pe_151_io_ve_out),
    .io_ho_out(bc_pe_151_io_ho_out),
    .io_res_out(bc_pe_151_io_res_out)
  );
  bc_pe bc_pe_152 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_152_clock),
    .reset(bc_pe_152_reset),
    .io_ho_input(bc_pe_152_io_ho_input),
    .io_ve_input(bc_pe_152_io_ve_input),
    .io_input_valid(bc_pe_152_io_input_valid),
    .io_iormac(bc_pe_152_io_iormac),
    .io_ve_out(bc_pe_152_io_ve_out),
    .io_ho_out(bc_pe_152_io_ho_out),
    .io_res_out(bc_pe_152_io_res_out)
  );
  bc_pe bc_pe_153 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_153_clock),
    .reset(bc_pe_153_reset),
    .io_ho_input(bc_pe_153_io_ho_input),
    .io_ve_input(bc_pe_153_io_ve_input),
    .io_input_valid(bc_pe_153_io_input_valid),
    .io_iormac(bc_pe_153_io_iormac),
    .io_ve_out(bc_pe_153_io_ve_out),
    .io_ho_out(bc_pe_153_io_ho_out),
    .io_res_out(bc_pe_153_io_res_out)
  );
  bc_pe bc_pe_154 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_154_clock),
    .reset(bc_pe_154_reset),
    .io_ho_input(bc_pe_154_io_ho_input),
    .io_ve_input(bc_pe_154_io_ve_input),
    .io_input_valid(bc_pe_154_io_input_valid),
    .io_iormac(bc_pe_154_io_iormac),
    .io_ve_out(bc_pe_154_io_ve_out),
    .io_ho_out(bc_pe_154_io_ho_out),
    .io_res_out(bc_pe_154_io_res_out)
  );
  bc_pe bc_pe_155 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_155_clock),
    .reset(bc_pe_155_reset),
    .io_ho_input(bc_pe_155_io_ho_input),
    .io_ve_input(bc_pe_155_io_ve_input),
    .io_input_valid(bc_pe_155_io_input_valid),
    .io_iormac(bc_pe_155_io_iormac),
    .io_ve_out(bc_pe_155_io_ve_out),
    .io_ho_out(bc_pe_155_io_ho_out),
    .io_res_out(bc_pe_155_io_res_out)
  );
  bc_pe bc_pe_156 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_156_clock),
    .reset(bc_pe_156_reset),
    .io_ho_input(bc_pe_156_io_ho_input),
    .io_ve_input(bc_pe_156_io_ve_input),
    .io_input_valid(bc_pe_156_io_input_valid),
    .io_iormac(bc_pe_156_io_iormac),
    .io_ve_out(bc_pe_156_io_ve_out),
    .io_ho_out(bc_pe_156_io_ho_out),
    .io_res_out(bc_pe_156_io_res_out)
  );
  bc_pe bc_pe_157 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_157_clock),
    .reset(bc_pe_157_reset),
    .io_ho_input(bc_pe_157_io_ho_input),
    .io_ve_input(bc_pe_157_io_ve_input),
    .io_input_valid(bc_pe_157_io_input_valid),
    .io_iormac(bc_pe_157_io_iormac),
    .io_ve_out(bc_pe_157_io_ve_out),
    .io_ho_out(bc_pe_157_io_ho_out),
    .io_res_out(bc_pe_157_io_res_out)
  );
  bc_pe bc_pe_158 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_158_clock),
    .reset(bc_pe_158_reset),
    .io_ho_input(bc_pe_158_io_ho_input),
    .io_ve_input(bc_pe_158_io_ve_input),
    .io_input_valid(bc_pe_158_io_input_valid),
    .io_iormac(bc_pe_158_io_iormac),
    .io_ve_out(bc_pe_158_io_ve_out),
    .io_ho_out(bc_pe_158_io_ho_out),
    .io_res_out(bc_pe_158_io_res_out)
  );
  bc_pe bc_pe_159 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_159_clock),
    .reset(bc_pe_159_reset),
    .io_ho_input(bc_pe_159_io_ho_input),
    .io_ve_input(bc_pe_159_io_ve_input),
    .io_input_valid(bc_pe_159_io_input_valid),
    .io_iormac(bc_pe_159_io_iormac),
    .io_ve_out(bc_pe_159_io_ve_out),
    .io_ho_out(bc_pe_159_io_ho_out),
    .io_res_out(bc_pe_159_io_res_out)
  );
  bc_pe bc_pe_160 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_160_clock),
    .reset(bc_pe_160_reset),
    .io_ho_input(bc_pe_160_io_ho_input),
    .io_ve_input(bc_pe_160_io_ve_input),
    .io_input_valid(bc_pe_160_io_input_valid),
    .io_iormac(bc_pe_160_io_iormac),
    .io_ve_out(bc_pe_160_io_ve_out),
    .io_ho_out(bc_pe_160_io_ho_out),
    .io_res_out(bc_pe_160_io_res_out)
  );
  bc_pe bc_pe_161 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_161_clock),
    .reset(bc_pe_161_reset),
    .io_ho_input(bc_pe_161_io_ho_input),
    .io_ve_input(bc_pe_161_io_ve_input),
    .io_input_valid(bc_pe_161_io_input_valid),
    .io_iormac(bc_pe_161_io_iormac),
    .io_ve_out(bc_pe_161_io_ve_out),
    .io_ho_out(bc_pe_161_io_ho_out),
    .io_res_out(bc_pe_161_io_res_out)
  );
  bc_pe bc_pe_162 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_162_clock),
    .reset(bc_pe_162_reset),
    .io_ho_input(bc_pe_162_io_ho_input),
    .io_ve_input(bc_pe_162_io_ve_input),
    .io_input_valid(bc_pe_162_io_input_valid),
    .io_iormac(bc_pe_162_io_iormac),
    .io_ve_out(bc_pe_162_io_ve_out),
    .io_ho_out(bc_pe_162_io_ho_out),
    .io_res_out(bc_pe_162_io_res_out)
  );
  bc_pe bc_pe_163 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_163_clock),
    .reset(bc_pe_163_reset),
    .io_ho_input(bc_pe_163_io_ho_input),
    .io_ve_input(bc_pe_163_io_ve_input),
    .io_input_valid(bc_pe_163_io_input_valid),
    .io_iormac(bc_pe_163_io_iormac),
    .io_ve_out(bc_pe_163_io_ve_out),
    .io_ho_out(bc_pe_163_io_ho_out),
    .io_res_out(bc_pe_163_io_res_out)
  );
  bc_pe bc_pe_164 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_164_clock),
    .reset(bc_pe_164_reset),
    .io_ho_input(bc_pe_164_io_ho_input),
    .io_ve_input(bc_pe_164_io_ve_input),
    .io_input_valid(bc_pe_164_io_input_valid),
    .io_iormac(bc_pe_164_io_iormac),
    .io_ve_out(bc_pe_164_io_ve_out),
    .io_ho_out(bc_pe_164_io_ho_out),
    .io_res_out(bc_pe_164_io_res_out)
  );
  bc_pe bc_pe_165 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_165_clock),
    .reset(bc_pe_165_reset),
    .io_ho_input(bc_pe_165_io_ho_input),
    .io_ve_input(bc_pe_165_io_ve_input),
    .io_input_valid(bc_pe_165_io_input_valid),
    .io_iormac(bc_pe_165_io_iormac),
    .io_ve_out(bc_pe_165_io_ve_out),
    .io_ho_out(bc_pe_165_io_ho_out),
    .io_res_out(bc_pe_165_io_res_out)
  );
  bc_pe bc_pe_166 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_166_clock),
    .reset(bc_pe_166_reset),
    .io_ho_input(bc_pe_166_io_ho_input),
    .io_ve_input(bc_pe_166_io_ve_input),
    .io_input_valid(bc_pe_166_io_input_valid),
    .io_iormac(bc_pe_166_io_iormac),
    .io_ve_out(bc_pe_166_io_ve_out),
    .io_ho_out(bc_pe_166_io_ho_out),
    .io_res_out(bc_pe_166_io_res_out)
  );
  bc_pe bc_pe_167 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_167_clock),
    .reset(bc_pe_167_reset),
    .io_ho_input(bc_pe_167_io_ho_input),
    .io_ve_input(bc_pe_167_io_ve_input),
    .io_input_valid(bc_pe_167_io_input_valid),
    .io_iormac(bc_pe_167_io_iormac),
    .io_ve_out(bc_pe_167_io_ve_out),
    .io_ho_out(bc_pe_167_io_ho_out),
    .io_res_out(bc_pe_167_io_res_out)
  );
  bc_pe bc_pe_168 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_168_clock),
    .reset(bc_pe_168_reset),
    .io_ho_input(bc_pe_168_io_ho_input),
    .io_ve_input(bc_pe_168_io_ve_input),
    .io_input_valid(bc_pe_168_io_input_valid),
    .io_iormac(bc_pe_168_io_iormac),
    .io_ve_out(bc_pe_168_io_ve_out),
    .io_ho_out(bc_pe_168_io_ho_out),
    .io_res_out(bc_pe_168_io_res_out)
  );
  bc_pe bc_pe_169 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_169_clock),
    .reset(bc_pe_169_reset),
    .io_ho_input(bc_pe_169_io_ho_input),
    .io_ve_input(bc_pe_169_io_ve_input),
    .io_input_valid(bc_pe_169_io_input_valid),
    .io_iormac(bc_pe_169_io_iormac),
    .io_ve_out(bc_pe_169_io_ve_out),
    .io_ho_out(bc_pe_169_io_ho_out),
    .io_res_out(bc_pe_169_io_res_out)
  );
  bc_pe bc_pe_170 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_170_clock),
    .reset(bc_pe_170_reset),
    .io_ho_input(bc_pe_170_io_ho_input),
    .io_ve_input(bc_pe_170_io_ve_input),
    .io_input_valid(bc_pe_170_io_input_valid),
    .io_iormac(bc_pe_170_io_iormac),
    .io_ve_out(bc_pe_170_io_ve_out),
    .io_ho_out(bc_pe_170_io_ho_out),
    .io_res_out(bc_pe_170_io_res_out)
  );
  bc_pe bc_pe_171 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_171_clock),
    .reset(bc_pe_171_reset),
    .io_ho_input(bc_pe_171_io_ho_input),
    .io_ve_input(bc_pe_171_io_ve_input),
    .io_input_valid(bc_pe_171_io_input_valid),
    .io_iormac(bc_pe_171_io_iormac),
    .io_ve_out(bc_pe_171_io_ve_out),
    .io_ho_out(bc_pe_171_io_ho_out),
    .io_res_out(bc_pe_171_io_res_out)
  );
  bc_pe bc_pe_172 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_172_clock),
    .reset(bc_pe_172_reset),
    .io_ho_input(bc_pe_172_io_ho_input),
    .io_ve_input(bc_pe_172_io_ve_input),
    .io_input_valid(bc_pe_172_io_input_valid),
    .io_iormac(bc_pe_172_io_iormac),
    .io_ve_out(bc_pe_172_io_ve_out),
    .io_ho_out(bc_pe_172_io_ho_out),
    .io_res_out(bc_pe_172_io_res_out)
  );
  bc_pe bc_pe_173 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_173_clock),
    .reset(bc_pe_173_reset),
    .io_ho_input(bc_pe_173_io_ho_input),
    .io_ve_input(bc_pe_173_io_ve_input),
    .io_input_valid(bc_pe_173_io_input_valid),
    .io_iormac(bc_pe_173_io_iormac),
    .io_ve_out(bc_pe_173_io_ve_out),
    .io_ho_out(bc_pe_173_io_ho_out),
    .io_res_out(bc_pe_173_io_res_out)
  );
  bc_pe bc_pe_174 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_174_clock),
    .reset(bc_pe_174_reset),
    .io_ho_input(bc_pe_174_io_ho_input),
    .io_ve_input(bc_pe_174_io_ve_input),
    .io_input_valid(bc_pe_174_io_input_valid),
    .io_iormac(bc_pe_174_io_iormac),
    .io_ve_out(bc_pe_174_io_ve_out),
    .io_ho_out(bc_pe_174_io_ho_out),
    .io_res_out(bc_pe_174_io_res_out)
  );
  bc_pe bc_pe_175 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_175_clock),
    .reset(bc_pe_175_reset),
    .io_ho_input(bc_pe_175_io_ho_input),
    .io_ve_input(bc_pe_175_io_ve_input),
    .io_input_valid(bc_pe_175_io_input_valid),
    .io_iormac(bc_pe_175_io_iormac),
    .io_ve_out(bc_pe_175_io_ve_out),
    .io_ho_out(bc_pe_175_io_ho_out),
    .io_res_out(bc_pe_175_io_res_out)
  );
  bc_pe bc_pe_176 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_176_clock),
    .reset(bc_pe_176_reset),
    .io_ho_input(bc_pe_176_io_ho_input),
    .io_ve_input(bc_pe_176_io_ve_input),
    .io_input_valid(bc_pe_176_io_input_valid),
    .io_iormac(bc_pe_176_io_iormac),
    .io_ve_out(bc_pe_176_io_ve_out),
    .io_ho_out(bc_pe_176_io_ho_out),
    .io_res_out(bc_pe_176_io_res_out)
  );
  bc_pe bc_pe_177 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_177_clock),
    .reset(bc_pe_177_reset),
    .io_ho_input(bc_pe_177_io_ho_input),
    .io_ve_input(bc_pe_177_io_ve_input),
    .io_input_valid(bc_pe_177_io_input_valid),
    .io_iormac(bc_pe_177_io_iormac),
    .io_ve_out(bc_pe_177_io_ve_out),
    .io_ho_out(bc_pe_177_io_ho_out),
    .io_res_out(bc_pe_177_io_res_out)
  );
  bc_pe bc_pe_178 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_178_clock),
    .reset(bc_pe_178_reset),
    .io_ho_input(bc_pe_178_io_ho_input),
    .io_ve_input(bc_pe_178_io_ve_input),
    .io_input_valid(bc_pe_178_io_input_valid),
    .io_iormac(bc_pe_178_io_iormac),
    .io_ve_out(bc_pe_178_io_ve_out),
    .io_ho_out(bc_pe_178_io_ho_out),
    .io_res_out(bc_pe_178_io_res_out)
  );
  bc_pe bc_pe_179 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_179_clock),
    .reset(bc_pe_179_reset),
    .io_ho_input(bc_pe_179_io_ho_input),
    .io_ve_input(bc_pe_179_io_ve_input),
    .io_input_valid(bc_pe_179_io_input_valid),
    .io_iormac(bc_pe_179_io_iormac),
    .io_ve_out(bc_pe_179_io_ve_out),
    .io_ho_out(bc_pe_179_io_ho_out),
    .io_res_out(bc_pe_179_io_res_out)
  );
  bc_pe bc_pe_180 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_180_clock),
    .reset(bc_pe_180_reset),
    .io_ho_input(bc_pe_180_io_ho_input),
    .io_ve_input(bc_pe_180_io_ve_input),
    .io_input_valid(bc_pe_180_io_input_valid),
    .io_iormac(bc_pe_180_io_iormac),
    .io_ve_out(bc_pe_180_io_ve_out),
    .io_ho_out(bc_pe_180_io_ho_out),
    .io_res_out(bc_pe_180_io_res_out)
  );
  bc_pe bc_pe_181 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_181_clock),
    .reset(bc_pe_181_reset),
    .io_ho_input(bc_pe_181_io_ho_input),
    .io_ve_input(bc_pe_181_io_ve_input),
    .io_input_valid(bc_pe_181_io_input_valid),
    .io_iormac(bc_pe_181_io_iormac),
    .io_ve_out(bc_pe_181_io_ve_out),
    .io_ho_out(bc_pe_181_io_ho_out),
    .io_res_out(bc_pe_181_io_res_out)
  );
  bc_pe bc_pe_182 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_182_clock),
    .reset(bc_pe_182_reset),
    .io_ho_input(bc_pe_182_io_ho_input),
    .io_ve_input(bc_pe_182_io_ve_input),
    .io_input_valid(bc_pe_182_io_input_valid),
    .io_iormac(bc_pe_182_io_iormac),
    .io_ve_out(bc_pe_182_io_ve_out),
    .io_ho_out(bc_pe_182_io_ho_out),
    .io_res_out(bc_pe_182_io_res_out)
  );
  bc_pe bc_pe_183 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_183_clock),
    .reset(bc_pe_183_reset),
    .io_ho_input(bc_pe_183_io_ho_input),
    .io_ve_input(bc_pe_183_io_ve_input),
    .io_input_valid(bc_pe_183_io_input_valid),
    .io_iormac(bc_pe_183_io_iormac),
    .io_ve_out(bc_pe_183_io_ve_out),
    .io_ho_out(bc_pe_183_io_ho_out),
    .io_res_out(bc_pe_183_io_res_out)
  );
  bc_pe bc_pe_184 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_184_clock),
    .reset(bc_pe_184_reset),
    .io_ho_input(bc_pe_184_io_ho_input),
    .io_ve_input(bc_pe_184_io_ve_input),
    .io_input_valid(bc_pe_184_io_input_valid),
    .io_iormac(bc_pe_184_io_iormac),
    .io_ve_out(bc_pe_184_io_ve_out),
    .io_ho_out(bc_pe_184_io_ho_out),
    .io_res_out(bc_pe_184_io_res_out)
  );
  bc_pe bc_pe_185 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_185_clock),
    .reset(bc_pe_185_reset),
    .io_ho_input(bc_pe_185_io_ho_input),
    .io_ve_input(bc_pe_185_io_ve_input),
    .io_input_valid(bc_pe_185_io_input_valid),
    .io_iormac(bc_pe_185_io_iormac),
    .io_ve_out(bc_pe_185_io_ve_out),
    .io_ho_out(bc_pe_185_io_ho_out),
    .io_res_out(bc_pe_185_io_res_out)
  );
  bc_pe bc_pe_186 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_186_clock),
    .reset(bc_pe_186_reset),
    .io_ho_input(bc_pe_186_io_ho_input),
    .io_ve_input(bc_pe_186_io_ve_input),
    .io_input_valid(bc_pe_186_io_input_valid),
    .io_iormac(bc_pe_186_io_iormac),
    .io_ve_out(bc_pe_186_io_ve_out),
    .io_ho_out(bc_pe_186_io_ho_out),
    .io_res_out(bc_pe_186_io_res_out)
  );
  bc_pe bc_pe_187 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_187_clock),
    .reset(bc_pe_187_reset),
    .io_ho_input(bc_pe_187_io_ho_input),
    .io_ve_input(bc_pe_187_io_ve_input),
    .io_input_valid(bc_pe_187_io_input_valid),
    .io_iormac(bc_pe_187_io_iormac),
    .io_ve_out(bc_pe_187_io_ve_out),
    .io_ho_out(bc_pe_187_io_ho_out),
    .io_res_out(bc_pe_187_io_res_out)
  );
  bc_pe bc_pe_188 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_188_clock),
    .reset(bc_pe_188_reset),
    .io_ho_input(bc_pe_188_io_ho_input),
    .io_ve_input(bc_pe_188_io_ve_input),
    .io_input_valid(bc_pe_188_io_input_valid),
    .io_iormac(bc_pe_188_io_iormac),
    .io_ve_out(bc_pe_188_io_ve_out),
    .io_ho_out(bc_pe_188_io_ho_out),
    .io_res_out(bc_pe_188_io_res_out)
  );
  bc_pe bc_pe_189 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_189_clock),
    .reset(bc_pe_189_reset),
    .io_ho_input(bc_pe_189_io_ho_input),
    .io_ve_input(bc_pe_189_io_ve_input),
    .io_input_valid(bc_pe_189_io_input_valid),
    .io_iormac(bc_pe_189_io_iormac),
    .io_ve_out(bc_pe_189_io_ve_out),
    .io_ho_out(bc_pe_189_io_ho_out),
    .io_res_out(bc_pe_189_io_res_out)
  );
  bc_pe bc_pe_190 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_190_clock),
    .reset(bc_pe_190_reset),
    .io_ho_input(bc_pe_190_io_ho_input),
    .io_ve_input(bc_pe_190_io_ve_input),
    .io_input_valid(bc_pe_190_io_input_valid),
    .io_iormac(bc_pe_190_io_iormac),
    .io_ve_out(bc_pe_190_io_ve_out),
    .io_ho_out(bc_pe_190_io_ho_out),
    .io_res_out(bc_pe_190_io_res_out)
  );
  bc_pe bc_pe_191 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_191_clock),
    .reset(bc_pe_191_reset),
    .io_ho_input(bc_pe_191_io_ho_input),
    .io_ve_input(bc_pe_191_io_ve_input),
    .io_input_valid(bc_pe_191_io_input_valid),
    .io_iormac(bc_pe_191_io_iormac),
    .io_ve_out(bc_pe_191_io_ve_out),
    .io_ho_out(bc_pe_191_io_ho_out),
    .io_res_out(bc_pe_191_io_res_out)
  );
  bc_pe bc_pe_192 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_192_clock),
    .reset(bc_pe_192_reset),
    .io_ho_input(bc_pe_192_io_ho_input),
    .io_ve_input(bc_pe_192_io_ve_input),
    .io_input_valid(bc_pe_192_io_input_valid),
    .io_iormac(bc_pe_192_io_iormac),
    .io_ve_out(bc_pe_192_io_ve_out),
    .io_ho_out(bc_pe_192_io_ho_out),
    .io_res_out(bc_pe_192_io_res_out)
  );
  bc_pe bc_pe_193 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_193_clock),
    .reset(bc_pe_193_reset),
    .io_ho_input(bc_pe_193_io_ho_input),
    .io_ve_input(bc_pe_193_io_ve_input),
    .io_input_valid(bc_pe_193_io_input_valid),
    .io_iormac(bc_pe_193_io_iormac),
    .io_ve_out(bc_pe_193_io_ve_out),
    .io_ho_out(bc_pe_193_io_ho_out),
    .io_res_out(bc_pe_193_io_res_out)
  );
  bc_pe bc_pe_194 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_194_clock),
    .reset(bc_pe_194_reset),
    .io_ho_input(bc_pe_194_io_ho_input),
    .io_ve_input(bc_pe_194_io_ve_input),
    .io_input_valid(bc_pe_194_io_input_valid),
    .io_iormac(bc_pe_194_io_iormac),
    .io_ve_out(bc_pe_194_io_ve_out),
    .io_ho_out(bc_pe_194_io_ho_out),
    .io_res_out(bc_pe_194_io_res_out)
  );
  bc_pe bc_pe_195 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_195_clock),
    .reset(bc_pe_195_reset),
    .io_ho_input(bc_pe_195_io_ho_input),
    .io_ve_input(bc_pe_195_io_ve_input),
    .io_input_valid(bc_pe_195_io_input_valid),
    .io_iormac(bc_pe_195_io_iormac),
    .io_ve_out(bc_pe_195_io_ve_out),
    .io_ho_out(bc_pe_195_io_ho_out),
    .io_res_out(bc_pe_195_io_res_out)
  );
  bc_pe bc_pe_196 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_196_clock),
    .reset(bc_pe_196_reset),
    .io_ho_input(bc_pe_196_io_ho_input),
    .io_ve_input(bc_pe_196_io_ve_input),
    .io_input_valid(bc_pe_196_io_input_valid),
    .io_iormac(bc_pe_196_io_iormac),
    .io_ve_out(bc_pe_196_io_ve_out),
    .io_ho_out(bc_pe_196_io_ho_out),
    .io_res_out(bc_pe_196_io_res_out)
  );
  bc_pe bc_pe_197 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_197_clock),
    .reset(bc_pe_197_reset),
    .io_ho_input(bc_pe_197_io_ho_input),
    .io_ve_input(bc_pe_197_io_ve_input),
    .io_input_valid(bc_pe_197_io_input_valid),
    .io_iormac(bc_pe_197_io_iormac),
    .io_ve_out(bc_pe_197_io_ve_out),
    .io_ho_out(bc_pe_197_io_ho_out),
    .io_res_out(bc_pe_197_io_res_out)
  );
  bc_pe bc_pe_198 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_198_clock),
    .reset(bc_pe_198_reset),
    .io_ho_input(bc_pe_198_io_ho_input),
    .io_ve_input(bc_pe_198_io_ve_input),
    .io_input_valid(bc_pe_198_io_input_valid),
    .io_iormac(bc_pe_198_io_iormac),
    .io_ve_out(bc_pe_198_io_ve_out),
    .io_ho_out(bc_pe_198_io_ho_out),
    .io_res_out(bc_pe_198_io_res_out)
  );
  bc_pe bc_pe_199 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_199_clock),
    .reset(bc_pe_199_reset),
    .io_ho_input(bc_pe_199_io_ho_input),
    .io_ve_input(bc_pe_199_io_ve_input),
    .io_input_valid(bc_pe_199_io_input_valid),
    .io_iormac(bc_pe_199_io_iormac),
    .io_ve_out(bc_pe_199_io_ve_out),
    .io_ho_out(bc_pe_199_io_ho_out),
    .io_res_out(bc_pe_199_io_res_out)
  );
  bc_pe bc_pe_200 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_200_clock),
    .reset(bc_pe_200_reset),
    .io_ho_input(bc_pe_200_io_ho_input),
    .io_ve_input(bc_pe_200_io_ve_input),
    .io_input_valid(bc_pe_200_io_input_valid),
    .io_iormac(bc_pe_200_io_iormac),
    .io_ve_out(bc_pe_200_io_ve_out),
    .io_ho_out(bc_pe_200_io_ho_out),
    .io_res_out(bc_pe_200_io_res_out)
  );
  bc_pe bc_pe_201 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_201_clock),
    .reset(bc_pe_201_reset),
    .io_ho_input(bc_pe_201_io_ho_input),
    .io_ve_input(bc_pe_201_io_ve_input),
    .io_input_valid(bc_pe_201_io_input_valid),
    .io_iormac(bc_pe_201_io_iormac),
    .io_ve_out(bc_pe_201_io_ve_out),
    .io_ho_out(bc_pe_201_io_ho_out),
    .io_res_out(bc_pe_201_io_res_out)
  );
  bc_pe bc_pe_202 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_202_clock),
    .reset(bc_pe_202_reset),
    .io_ho_input(bc_pe_202_io_ho_input),
    .io_ve_input(bc_pe_202_io_ve_input),
    .io_input_valid(bc_pe_202_io_input_valid),
    .io_iormac(bc_pe_202_io_iormac),
    .io_ve_out(bc_pe_202_io_ve_out),
    .io_ho_out(bc_pe_202_io_ho_out),
    .io_res_out(bc_pe_202_io_res_out)
  );
  bc_pe bc_pe_203 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_203_clock),
    .reset(bc_pe_203_reset),
    .io_ho_input(bc_pe_203_io_ho_input),
    .io_ve_input(bc_pe_203_io_ve_input),
    .io_input_valid(bc_pe_203_io_input_valid),
    .io_iormac(bc_pe_203_io_iormac),
    .io_ve_out(bc_pe_203_io_ve_out),
    .io_ho_out(bc_pe_203_io_ho_out),
    .io_res_out(bc_pe_203_io_res_out)
  );
  bc_pe bc_pe_204 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_204_clock),
    .reset(bc_pe_204_reset),
    .io_ho_input(bc_pe_204_io_ho_input),
    .io_ve_input(bc_pe_204_io_ve_input),
    .io_input_valid(bc_pe_204_io_input_valid),
    .io_iormac(bc_pe_204_io_iormac),
    .io_ve_out(bc_pe_204_io_ve_out),
    .io_ho_out(bc_pe_204_io_ho_out),
    .io_res_out(bc_pe_204_io_res_out)
  );
  bc_pe bc_pe_205 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_205_clock),
    .reset(bc_pe_205_reset),
    .io_ho_input(bc_pe_205_io_ho_input),
    .io_ve_input(bc_pe_205_io_ve_input),
    .io_input_valid(bc_pe_205_io_input_valid),
    .io_iormac(bc_pe_205_io_iormac),
    .io_ve_out(bc_pe_205_io_ve_out),
    .io_ho_out(bc_pe_205_io_ho_out),
    .io_res_out(bc_pe_205_io_res_out)
  );
  bc_pe bc_pe_206 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_206_clock),
    .reset(bc_pe_206_reset),
    .io_ho_input(bc_pe_206_io_ho_input),
    .io_ve_input(bc_pe_206_io_ve_input),
    .io_input_valid(bc_pe_206_io_input_valid),
    .io_iormac(bc_pe_206_io_iormac),
    .io_ve_out(bc_pe_206_io_ve_out),
    .io_ho_out(bc_pe_206_io_ho_out),
    .io_res_out(bc_pe_206_io_res_out)
  );
  bc_pe bc_pe_207 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_207_clock),
    .reset(bc_pe_207_reset),
    .io_ho_input(bc_pe_207_io_ho_input),
    .io_ve_input(bc_pe_207_io_ve_input),
    .io_input_valid(bc_pe_207_io_input_valid),
    .io_iormac(bc_pe_207_io_iormac),
    .io_ve_out(bc_pe_207_io_ve_out),
    .io_ho_out(bc_pe_207_io_ho_out),
    .io_res_out(bc_pe_207_io_res_out)
  );
  bc_pe bc_pe_208 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_208_clock),
    .reset(bc_pe_208_reset),
    .io_ho_input(bc_pe_208_io_ho_input),
    .io_ve_input(bc_pe_208_io_ve_input),
    .io_input_valid(bc_pe_208_io_input_valid),
    .io_iormac(bc_pe_208_io_iormac),
    .io_ve_out(bc_pe_208_io_ve_out),
    .io_ho_out(bc_pe_208_io_ho_out),
    .io_res_out(bc_pe_208_io_res_out)
  );
  bc_pe bc_pe_209 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_209_clock),
    .reset(bc_pe_209_reset),
    .io_ho_input(bc_pe_209_io_ho_input),
    .io_ve_input(bc_pe_209_io_ve_input),
    .io_input_valid(bc_pe_209_io_input_valid),
    .io_iormac(bc_pe_209_io_iormac),
    .io_ve_out(bc_pe_209_io_ve_out),
    .io_ho_out(bc_pe_209_io_ho_out),
    .io_res_out(bc_pe_209_io_res_out)
  );
  bc_pe bc_pe_210 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_210_clock),
    .reset(bc_pe_210_reset),
    .io_ho_input(bc_pe_210_io_ho_input),
    .io_ve_input(bc_pe_210_io_ve_input),
    .io_input_valid(bc_pe_210_io_input_valid),
    .io_iormac(bc_pe_210_io_iormac),
    .io_ve_out(bc_pe_210_io_ve_out),
    .io_ho_out(bc_pe_210_io_ho_out),
    .io_res_out(bc_pe_210_io_res_out)
  );
  bc_pe bc_pe_211 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_211_clock),
    .reset(bc_pe_211_reset),
    .io_ho_input(bc_pe_211_io_ho_input),
    .io_ve_input(bc_pe_211_io_ve_input),
    .io_input_valid(bc_pe_211_io_input_valid),
    .io_iormac(bc_pe_211_io_iormac),
    .io_ve_out(bc_pe_211_io_ve_out),
    .io_ho_out(bc_pe_211_io_ho_out),
    .io_res_out(bc_pe_211_io_res_out)
  );
  bc_pe bc_pe_212 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_212_clock),
    .reset(bc_pe_212_reset),
    .io_ho_input(bc_pe_212_io_ho_input),
    .io_ve_input(bc_pe_212_io_ve_input),
    .io_input_valid(bc_pe_212_io_input_valid),
    .io_iormac(bc_pe_212_io_iormac),
    .io_ve_out(bc_pe_212_io_ve_out),
    .io_ho_out(bc_pe_212_io_ho_out),
    .io_res_out(bc_pe_212_io_res_out)
  );
  bc_pe bc_pe_213 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_213_clock),
    .reset(bc_pe_213_reset),
    .io_ho_input(bc_pe_213_io_ho_input),
    .io_ve_input(bc_pe_213_io_ve_input),
    .io_input_valid(bc_pe_213_io_input_valid),
    .io_iormac(bc_pe_213_io_iormac),
    .io_ve_out(bc_pe_213_io_ve_out),
    .io_ho_out(bc_pe_213_io_ho_out),
    .io_res_out(bc_pe_213_io_res_out)
  );
  bc_pe bc_pe_214 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_214_clock),
    .reset(bc_pe_214_reset),
    .io_ho_input(bc_pe_214_io_ho_input),
    .io_ve_input(bc_pe_214_io_ve_input),
    .io_input_valid(bc_pe_214_io_input_valid),
    .io_iormac(bc_pe_214_io_iormac),
    .io_ve_out(bc_pe_214_io_ve_out),
    .io_ho_out(bc_pe_214_io_ho_out),
    .io_res_out(bc_pe_214_io_res_out)
  );
  bc_pe bc_pe_215 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_215_clock),
    .reset(bc_pe_215_reset),
    .io_ho_input(bc_pe_215_io_ho_input),
    .io_ve_input(bc_pe_215_io_ve_input),
    .io_input_valid(bc_pe_215_io_input_valid),
    .io_iormac(bc_pe_215_io_iormac),
    .io_ve_out(bc_pe_215_io_ve_out),
    .io_ho_out(bc_pe_215_io_ho_out),
    .io_res_out(bc_pe_215_io_res_out)
  );
  bc_pe bc_pe_216 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_216_clock),
    .reset(bc_pe_216_reset),
    .io_ho_input(bc_pe_216_io_ho_input),
    .io_ve_input(bc_pe_216_io_ve_input),
    .io_input_valid(bc_pe_216_io_input_valid),
    .io_iormac(bc_pe_216_io_iormac),
    .io_ve_out(bc_pe_216_io_ve_out),
    .io_ho_out(bc_pe_216_io_ho_out),
    .io_res_out(bc_pe_216_io_res_out)
  );
  bc_pe bc_pe_217 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_217_clock),
    .reset(bc_pe_217_reset),
    .io_ho_input(bc_pe_217_io_ho_input),
    .io_ve_input(bc_pe_217_io_ve_input),
    .io_input_valid(bc_pe_217_io_input_valid),
    .io_iormac(bc_pe_217_io_iormac),
    .io_ve_out(bc_pe_217_io_ve_out),
    .io_ho_out(bc_pe_217_io_ho_out),
    .io_res_out(bc_pe_217_io_res_out)
  );
  bc_pe bc_pe_218 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_218_clock),
    .reset(bc_pe_218_reset),
    .io_ho_input(bc_pe_218_io_ho_input),
    .io_ve_input(bc_pe_218_io_ve_input),
    .io_input_valid(bc_pe_218_io_input_valid),
    .io_iormac(bc_pe_218_io_iormac),
    .io_ve_out(bc_pe_218_io_ve_out),
    .io_ho_out(bc_pe_218_io_ho_out),
    .io_res_out(bc_pe_218_io_res_out)
  );
  bc_pe bc_pe_219 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_219_clock),
    .reset(bc_pe_219_reset),
    .io_ho_input(bc_pe_219_io_ho_input),
    .io_ve_input(bc_pe_219_io_ve_input),
    .io_input_valid(bc_pe_219_io_input_valid),
    .io_iormac(bc_pe_219_io_iormac),
    .io_ve_out(bc_pe_219_io_ve_out),
    .io_ho_out(bc_pe_219_io_ho_out),
    .io_res_out(bc_pe_219_io_res_out)
  );
  bc_pe bc_pe_220 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_220_clock),
    .reset(bc_pe_220_reset),
    .io_ho_input(bc_pe_220_io_ho_input),
    .io_ve_input(bc_pe_220_io_ve_input),
    .io_input_valid(bc_pe_220_io_input_valid),
    .io_iormac(bc_pe_220_io_iormac),
    .io_ve_out(bc_pe_220_io_ve_out),
    .io_ho_out(bc_pe_220_io_ho_out),
    .io_res_out(bc_pe_220_io_res_out)
  );
  bc_pe bc_pe_221 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_221_clock),
    .reset(bc_pe_221_reset),
    .io_ho_input(bc_pe_221_io_ho_input),
    .io_ve_input(bc_pe_221_io_ve_input),
    .io_input_valid(bc_pe_221_io_input_valid),
    .io_iormac(bc_pe_221_io_iormac),
    .io_ve_out(bc_pe_221_io_ve_out),
    .io_ho_out(bc_pe_221_io_ho_out),
    .io_res_out(bc_pe_221_io_res_out)
  );
  bc_pe bc_pe_222 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_222_clock),
    .reset(bc_pe_222_reset),
    .io_ho_input(bc_pe_222_io_ho_input),
    .io_ve_input(bc_pe_222_io_ve_input),
    .io_input_valid(bc_pe_222_io_input_valid),
    .io_iormac(bc_pe_222_io_iormac),
    .io_ve_out(bc_pe_222_io_ve_out),
    .io_ho_out(bc_pe_222_io_ho_out),
    .io_res_out(bc_pe_222_io_res_out)
  );
  bc_pe bc_pe_223 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_223_clock),
    .reset(bc_pe_223_reset),
    .io_ho_input(bc_pe_223_io_ho_input),
    .io_ve_input(bc_pe_223_io_ve_input),
    .io_input_valid(bc_pe_223_io_input_valid),
    .io_iormac(bc_pe_223_io_iormac),
    .io_ve_out(bc_pe_223_io_ve_out),
    .io_ho_out(bc_pe_223_io_ho_out),
    .io_res_out(bc_pe_223_io_res_out)
  );
  bc_pe bc_pe_224 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_224_clock),
    .reset(bc_pe_224_reset),
    .io_ho_input(bc_pe_224_io_ho_input),
    .io_ve_input(bc_pe_224_io_ve_input),
    .io_input_valid(bc_pe_224_io_input_valid),
    .io_iormac(bc_pe_224_io_iormac),
    .io_ve_out(bc_pe_224_io_ve_out),
    .io_ho_out(bc_pe_224_io_ho_out),
    .io_res_out(bc_pe_224_io_res_out)
  );
  bc_pe bc_pe_225 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_225_clock),
    .reset(bc_pe_225_reset),
    .io_ho_input(bc_pe_225_io_ho_input),
    .io_ve_input(bc_pe_225_io_ve_input),
    .io_input_valid(bc_pe_225_io_input_valid),
    .io_iormac(bc_pe_225_io_iormac),
    .io_ve_out(bc_pe_225_io_ve_out),
    .io_ho_out(bc_pe_225_io_ho_out),
    .io_res_out(bc_pe_225_io_res_out)
  );
  bc_pe bc_pe_226 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_226_clock),
    .reset(bc_pe_226_reset),
    .io_ho_input(bc_pe_226_io_ho_input),
    .io_ve_input(bc_pe_226_io_ve_input),
    .io_input_valid(bc_pe_226_io_input_valid),
    .io_iormac(bc_pe_226_io_iormac),
    .io_ve_out(bc_pe_226_io_ve_out),
    .io_ho_out(bc_pe_226_io_ho_out),
    .io_res_out(bc_pe_226_io_res_out)
  );
  bc_pe bc_pe_227 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_227_clock),
    .reset(bc_pe_227_reset),
    .io_ho_input(bc_pe_227_io_ho_input),
    .io_ve_input(bc_pe_227_io_ve_input),
    .io_input_valid(bc_pe_227_io_input_valid),
    .io_iormac(bc_pe_227_io_iormac),
    .io_ve_out(bc_pe_227_io_ve_out),
    .io_ho_out(bc_pe_227_io_ho_out),
    .io_res_out(bc_pe_227_io_res_out)
  );
  bc_pe bc_pe_228 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_228_clock),
    .reset(bc_pe_228_reset),
    .io_ho_input(bc_pe_228_io_ho_input),
    .io_ve_input(bc_pe_228_io_ve_input),
    .io_input_valid(bc_pe_228_io_input_valid),
    .io_iormac(bc_pe_228_io_iormac),
    .io_ve_out(bc_pe_228_io_ve_out),
    .io_ho_out(bc_pe_228_io_ho_out),
    .io_res_out(bc_pe_228_io_res_out)
  );
  bc_pe bc_pe_229 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_229_clock),
    .reset(bc_pe_229_reset),
    .io_ho_input(bc_pe_229_io_ho_input),
    .io_ve_input(bc_pe_229_io_ve_input),
    .io_input_valid(bc_pe_229_io_input_valid),
    .io_iormac(bc_pe_229_io_iormac),
    .io_ve_out(bc_pe_229_io_ve_out),
    .io_ho_out(bc_pe_229_io_ho_out),
    .io_res_out(bc_pe_229_io_res_out)
  );
  bc_pe bc_pe_230 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_230_clock),
    .reset(bc_pe_230_reset),
    .io_ho_input(bc_pe_230_io_ho_input),
    .io_ve_input(bc_pe_230_io_ve_input),
    .io_input_valid(bc_pe_230_io_input_valid),
    .io_iormac(bc_pe_230_io_iormac),
    .io_ve_out(bc_pe_230_io_ve_out),
    .io_ho_out(bc_pe_230_io_ho_out),
    .io_res_out(bc_pe_230_io_res_out)
  );
  bc_pe bc_pe_231 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_231_clock),
    .reset(bc_pe_231_reset),
    .io_ho_input(bc_pe_231_io_ho_input),
    .io_ve_input(bc_pe_231_io_ve_input),
    .io_input_valid(bc_pe_231_io_input_valid),
    .io_iormac(bc_pe_231_io_iormac),
    .io_ve_out(bc_pe_231_io_ve_out),
    .io_ho_out(bc_pe_231_io_ho_out),
    .io_res_out(bc_pe_231_io_res_out)
  );
  bc_pe bc_pe_232 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_232_clock),
    .reset(bc_pe_232_reset),
    .io_ho_input(bc_pe_232_io_ho_input),
    .io_ve_input(bc_pe_232_io_ve_input),
    .io_input_valid(bc_pe_232_io_input_valid),
    .io_iormac(bc_pe_232_io_iormac),
    .io_ve_out(bc_pe_232_io_ve_out),
    .io_ho_out(bc_pe_232_io_ho_out),
    .io_res_out(bc_pe_232_io_res_out)
  );
  bc_pe bc_pe_233 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_233_clock),
    .reset(bc_pe_233_reset),
    .io_ho_input(bc_pe_233_io_ho_input),
    .io_ve_input(bc_pe_233_io_ve_input),
    .io_input_valid(bc_pe_233_io_input_valid),
    .io_iormac(bc_pe_233_io_iormac),
    .io_ve_out(bc_pe_233_io_ve_out),
    .io_ho_out(bc_pe_233_io_ho_out),
    .io_res_out(bc_pe_233_io_res_out)
  );
  bc_pe bc_pe_234 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_234_clock),
    .reset(bc_pe_234_reset),
    .io_ho_input(bc_pe_234_io_ho_input),
    .io_ve_input(bc_pe_234_io_ve_input),
    .io_input_valid(bc_pe_234_io_input_valid),
    .io_iormac(bc_pe_234_io_iormac),
    .io_ve_out(bc_pe_234_io_ve_out),
    .io_ho_out(bc_pe_234_io_ho_out),
    .io_res_out(bc_pe_234_io_res_out)
  );
  bc_pe bc_pe_235 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_235_clock),
    .reset(bc_pe_235_reset),
    .io_ho_input(bc_pe_235_io_ho_input),
    .io_ve_input(bc_pe_235_io_ve_input),
    .io_input_valid(bc_pe_235_io_input_valid),
    .io_iormac(bc_pe_235_io_iormac),
    .io_ve_out(bc_pe_235_io_ve_out),
    .io_ho_out(bc_pe_235_io_ho_out),
    .io_res_out(bc_pe_235_io_res_out)
  );
  bc_pe bc_pe_236 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_236_clock),
    .reset(bc_pe_236_reset),
    .io_ho_input(bc_pe_236_io_ho_input),
    .io_ve_input(bc_pe_236_io_ve_input),
    .io_input_valid(bc_pe_236_io_input_valid),
    .io_iormac(bc_pe_236_io_iormac),
    .io_ve_out(bc_pe_236_io_ve_out),
    .io_ho_out(bc_pe_236_io_ho_out),
    .io_res_out(bc_pe_236_io_res_out)
  );
  bc_pe bc_pe_237 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_237_clock),
    .reset(bc_pe_237_reset),
    .io_ho_input(bc_pe_237_io_ho_input),
    .io_ve_input(bc_pe_237_io_ve_input),
    .io_input_valid(bc_pe_237_io_input_valid),
    .io_iormac(bc_pe_237_io_iormac),
    .io_ve_out(bc_pe_237_io_ve_out),
    .io_ho_out(bc_pe_237_io_ho_out),
    .io_res_out(bc_pe_237_io_res_out)
  );
  bc_pe bc_pe_238 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_238_clock),
    .reset(bc_pe_238_reset),
    .io_ho_input(bc_pe_238_io_ho_input),
    .io_ve_input(bc_pe_238_io_ve_input),
    .io_input_valid(bc_pe_238_io_input_valid),
    .io_iormac(bc_pe_238_io_iormac),
    .io_ve_out(bc_pe_238_io_ve_out),
    .io_ho_out(bc_pe_238_io_ho_out),
    .io_res_out(bc_pe_238_io_res_out)
  );
  bc_pe bc_pe_239 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_239_clock),
    .reset(bc_pe_239_reset),
    .io_ho_input(bc_pe_239_io_ho_input),
    .io_ve_input(bc_pe_239_io_ve_input),
    .io_input_valid(bc_pe_239_io_input_valid),
    .io_iormac(bc_pe_239_io_iormac),
    .io_ve_out(bc_pe_239_io_ve_out),
    .io_ho_out(bc_pe_239_io_ho_out),
    .io_res_out(bc_pe_239_io_res_out)
  );
  bc_pe bc_pe_240 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_240_clock),
    .reset(bc_pe_240_reset),
    .io_ho_input(bc_pe_240_io_ho_input),
    .io_ve_input(bc_pe_240_io_ve_input),
    .io_input_valid(bc_pe_240_io_input_valid),
    .io_iormac(bc_pe_240_io_iormac),
    .io_ve_out(bc_pe_240_io_ve_out),
    .io_ho_out(bc_pe_240_io_ho_out),
    .io_res_out(bc_pe_240_io_res_out)
  );
  bc_pe bc_pe_241 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_241_clock),
    .reset(bc_pe_241_reset),
    .io_ho_input(bc_pe_241_io_ho_input),
    .io_ve_input(bc_pe_241_io_ve_input),
    .io_input_valid(bc_pe_241_io_input_valid),
    .io_iormac(bc_pe_241_io_iormac),
    .io_ve_out(bc_pe_241_io_ve_out),
    .io_ho_out(bc_pe_241_io_ho_out),
    .io_res_out(bc_pe_241_io_res_out)
  );
  bc_pe bc_pe_242 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_242_clock),
    .reset(bc_pe_242_reset),
    .io_ho_input(bc_pe_242_io_ho_input),
    .io_ve_input(bc_pe_242_io_ve_input),
    .io_input_valid(bc_pe_242_io_input_valid),
    .io_iormac(bc_pe_242_io_iormac),
    .io_ve_out(bc_pe_242_io_ve_out),
    .io_ho_out(bc_pe_242_io_ho_out),
    .io_res_out(bc_pe_242_io_res_out)
  );
  bc_pe bc_pe_243 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_243_clock),
    .reset(bc_pe_243_reset),
    .io_ho_input(bc_pe_243_io_ho_input),
    .io_ve_input(bc_pe_243_io_ve_input),
    .io_input_valid(bc_pe_243_io_input_valid),
    .io_iormac(bc_pe_243_io_iormac),
    .io_ve_out(bc_pe_243_io_ve_out),
    .io_ho_out(bc_pe_243_io_ho_out),
    .io_res_out(bc_pe_243_io_res_out)
  );
  bc_pe bc_pe_244 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_244_clock),
    .reset(bc_pe_244_reset),
    .io_ho_input(bc_pe_244_io_ho_input),
    .io_ve_input(bc_pe_244_io_ve_input),
    .io_input_valid(bc_pe_244_io_input_valid),
    .io_iormac(bc_pe_244_io_iormac),
    .io_ve_out(bc_pe_244_io_ve_out),
    .io_ho_out(bc_pe_244_io_ho_out),
    .io_res_out(bc_pe_244_io_res_out)
  );
  bc_pe bc_pe_245 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_245_clock),
    .reset(bc_pe_245_reset),
    .io_ho_input(bc_pe_245_io_ho_input),
    .io_ve_input(bc_pe_245_io_ve_input),
    .io_input_valid(bc_pe_245_io_input_valid),
    .io_iormac(bc_pe_245_io_iormac),
    .io_ve_out(bc_pe_245_io_ve_out),
    .io_ho_out(bc_pe_245_io_ho_out),
    .io_res_out(bc_pe_245_io_res_out)
  );
  bc_pe bc_pe_246 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_246_clock),
    .reset(bc_pe_246_reset),
    .io_ho_input(bc_pe_246_io_ho_input),
    .io_ve_input(bc_pe_246_io_ve_input),
    .io_input_valid(bc_pe_246_io_input_valid),
    .io_iormac(bc_pe_246_io_iormac),
    .io_ve_out(bc_pe_246_io_ve_out),
    .io_ho_out(bc_pe_246_io_ho_out),
    .io_res_out(bc_pe_246_io_res_out)
  );
  bc_pe bc_pe_247 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_247_clock),
    .reset(bc_pe_247_reset),
    .io_ho_input(bc_pe_247_io_ho_input),
    .io_ve_input(bc_pe_247_io_ve_input),
    .io_input_valid(bc_pe_247_io_input_valid),
    .io_iormac(bc_pe_247_io_iormac),
    .io_ve_out(bc_pe_247_io_ve_out),
    .io_ho_out(bc_pe_247_io_ho_out),
    .io_res_out(bc_pe_247_io_res_out)
  );
  bc_pe bc_pe_248 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_248_clock),
    .reset(bc_pe_248_reset),
    .io_ho_input(bc_pe_248_io_ho_input),
    .io_ve_input(bc_pe_248_io_ve_input),
    .io_input_valid(bc_pe_248_io_input_valid),
    .io_iormac(bc_pe_248_io_iormac),
    .io_ve_out(bc_pe_248_io_ve_out),
    .io_ho_out(bc_pe_248_io_ho_out),
    .io_res_out(bc_pe_248_io_res_out)
  );
  bc_pe bc_pe_249 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_249_clock),
    .reset(bc_pe_249_reset),
    .io_ho_input(bc_pe_249_io_ho_input),
    .io_ve_input(bc_pe_249_io_ve_input),
    .io_input_valid(bc_pe_249_io_input_valid),
    .io_iormac(bc_pe_249_io_iormac),
    .io_ve_out(bc_pe_249_io_ve_out),
    .io_ho_out(bc_pe_249_io_ho_out),
    .io_res_out(bc_pe_249_io_res_out)
  );
  bc_pe bc_pe_250 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_250_clock),
    .reset(bc_pe_250_reset),
    .io_ho_input(bc_pe_250_io_ho_input),
    .io_ve_input(bc_pe_250_io_ve_input),
    .io_input_valid(bc_pe_250_io_input_valid),
    .io_iormac(bc_pe_250_io_iormac),
    .io_ve_out(bc_pe_250_io_ve_out),
    .io_ho_out(bc_pe_250_io_ho_out),
    .io_res_out(bc_pe_250_io_res_out)
  );
  bc_pe bc_pe_251 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_251_clock),
    .reset(bc_pe_251_reset),
    .io_ho_input(bc_pe_251_io_ho_input),
    .io_ve_input(bc_pe_251_io_ve_input),
    .io_input_valid(bc_pe_251_io_input_valid),
    .io_iormac(bc_pe_251_io_iormac),
    .io_ve_out(bc_pe_251_io_ve_out),
    .io_ho_out(bc_pe_251_io_ho_out),
    .io_res_out(bc_pe_251_io_res_out)
  );
  bc_pe bc_pe_252 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_252_clock),
    .reset(bc_pe_252_reset),
    .io_ho_input(bc_pe_252_io_ho_input),
    .io_ve_input(bc_pe_252_io_ve_input),
    .io_input_valid(bc_pe_252_io_input_valid),
    .io_iormac(bc_pe_252_io_iormac),
    .io_ve_out(bc_pe_252_io_ve_out),
    .io_ho_out(bc_pe_252_io_ho_out),
    .io_res_out(bc_pe_252_io_res_out)
  );
  bc_pe bc_pe_253 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_253_clock),
    .reset(bc_pe_253_reset),
    .io_ho_input(bc_pe_253_io_ho_input),
    .io_ve_input(bc_pe_253_io_ve_input),
    .io_input_valid(bc_pe_253_io_input_valid),
    .io_iormac(bc_pe_253_io_iormac),
    .io_ve_out(bc_pe_253_io_ve_out),
    .io_ho_out(bc_pe_253_io_ho_out),
    .io_res_out(bc_pe_253_io_res_out)
  );
  bc_pe bc_pe_254 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_254_clock),
    .reset(bc_pe_254_reset),
    .io_ho_input(bc_pe_254_io_ho_input),
    .io_ve_input(bc_pe_254_io_ve_input),
    .io_input_valid(bc_pe_254_io_input_valid),
    .io_iormac(bc_pe_254_io_iormac),
    .io_ve_out(bc_pe_254_io_ve_out),
    .io_ho_out(bc_pe_254_io_ho_out),
    .io_res_out(bc_pe_254_io_res_out)
  );
  bc_pe bc_pe_255 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_255_clock),
    .reset(bc_pe_255_reset),
    .io_ho_input(bc_pe_255_io_ho_input),
    .io_ve_input(bc_pe_255_io_ve_input),
    .io_input_valid(bc_pe_255_io_input_valid),
    .io_iormac(bc_pe_255_io_iormac),
    .io_ve_out(bc_pe_255_io_ve_out),
    .io_ho_out(bc_pe_255_io_ho_out),
    .io_res_out(bc_pe_255_io_res_out)
  );
  bc_pe bc_pe_256 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_256_clock),
    .reset(bc_pe_256_reset),
    .io_ho_input(bc_pe_256_io_ho_input),
    .io_ve_input(bc_pe_256_io_ve_input),
    .io_input_valid(bc_pe_256_io_input_valid),
    .io_iormac(bc_pe_256_io_iormac),
    .io_ve_out(bc_pe_256_io_ve_out),
    .io_ho_out(bc_pe_256_io_ho_out),
    .io_res_out(bc_pe_256_io_res_out)
  );
  bc_pe bc_pe_257 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_257_clock),
    .reset(bc_pe_257_reset),
    .io_ho_input(bc_pe_257_io_ho_input),
    .io_ve_input(bc_pe_257_io_ve_input),
    .io_input_valid(bc_pe_257_io_input_valid),
    .io_iormac(bc_pe_257_io_iormac),
    .io_ve_out(bc_pe_257_io_ve_out),
    .io_ho_out(bc_pe_257_io_ho_out),
    .io_res_out(bc_pe_257_io_res_out)
  );
  bc_pe bc_pe_258 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_258_clock),
    .reset(bc_pe_258_reset),
    .io_ho_input(bc_pe_258_io_ho_input),
    .io_ve_input(bc_pe_258_io_ve_input),
    .io_input_valid(bc_pe_258_io_input_valid),
    .io_iormac(bc_pe_258_io_iormac),
    .io_ve_out(bc_pe_258_io_ve_out),
    .io_ho_out(bc_pe_258_io_ho_out),
    .io_res_out(bc_pe_258_io_res_out)
  );
  bc_pe bc_pe_259 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_259_clock),
    .reset(bc_pe_259_reset),
    .io_ho_input(bc_pe_259_io_ho_input),
    .io_ve_input(bc_pe_259_io_ve_input),
    .io_input_valid(bc_pe_259_io_input_valid),
    .io_iormac(bc_pe_259_io_iormac),
    .io_ve_out(bc_pe_259_io_ve_out),
    .io_ho_out(bc_pe_259_io_ho_out),
    .io_res_out(bc_pe_259_io_res_out)
  );
  bc_pe bc_pe_260 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_260_clock),
    .reset(bc_pe_260_reset),
    .io_ho_input(bc_pe_260_io_ho_input),
    .io_ve_input(bc_pe_260_io_ve_input),
    .io_input_valid(bc_pe_260_io_input_valid),
    .io_iormac(bc_pe_260_io_iormac),
    .io_ve_out(bc_pe_260_io_ve_out),
    .io_ho_out(bc_pe_260_io_ho_out),
    .io_res_out(bc_pe_260_io_res_out)
  );
  bc_pe bc_pe_261 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_261_clock),
    .reset(bc_pe_261_reset),
    .io_ho_input(bc_pe_261_io_ho_input),
    .io_ve_input(bc_pe_261_io_ve_input),
    .io_input_valid(bc_pe_261_io_input_valid),
    .io_iormac(bc_pe_261_io_iormac),
    .io_ve_out(bc_pe_261_io_ve_out),
    .io_ho_out(bc_pe_261_io_ho_out),
    .io_res_out(bc_pe_261_io_res_out)
  );
  bc_pe bc_pe_262 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_262_clock),
    .reset(bc_pe_262_reset),
    .io_ho_input(bc_pe_262_io_ho_input),
    .io_ve_input(bc_pe_262_io_ve_input),
    .io_input_valid(bc_pe_262_io_input_valid),
    .io_iormac(bc_pe_262_io_iormac),
    .io_ve_out(bc_pe_262_io_ve_out),
    .io_ho_out(bc_pe_262_io_ho_out),
    .io_res_out(bc_pe_262_io_res_out)
  );
  bc_pe bc_pe_263 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_263_clock),
    .reset(bc_pe_263_reset),
    .io_ho_input(bc_pe_263_io_ho_input),
    .io_ve_input(bc_pe_263_io_ve_input),
    .io_input_valid(bc_pe_263_io_input_valid),
    .io_iormac(bc_pe_263_io_iormac),
    .io_ve_out(bc_pe_263_io_ve_out),
    .io_ho_out(bc_pe_263_io_ho_out),
    .io_res_out(bc_pe_263_io_res_out)
  );
  bc_pe bc_pe_264 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_264_clock),
    .reset(bc_pe_264_reset),
    .io_ho_input(bc_pe_264_io_ho_input),
    .io_ve_input(bc_pe_264_io_ve_input),
    .io_input_valid(bc_pe_264_io_input_valid),
    .io_iormac(bc_pe_264_io_iormac),
    .io_ve_out(bc_pe_264_io_ve_out),
    .io_ho_out(bc_pe_264_io_ho_out),
    .io_res_out(bc_pe_264_io_res_out)
  );
  bc_pe bc_pe_265 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_265_clock),
    .reset(bc_pe_265_reset),
    .io_ho_input(bc_pe_265_io_ho_input),
    .io_ve_input(bc_pe_265_io_ve_input),
    .io_input_valid(bc_pe_265_io_input_valid),
    .io_iormac(bc_pe_265_io_iormac),
    .io_ve_out(bc_pe_265_io_ve_out),
    .io_ho_out(bc_pe_265_io_ho_out),
    .io_res_out(bc_pe_265_io_res_out)
  );
  bc_pe bc_pe_266 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_266_clock),
    .reset(bc_pe_266_reset),
    .io_ho_input(bc_pe_266_io_ho_input),
    .io_ve_input(bc_pe_266_io_ve_input),
    .io_input_valid(bc_pe_266_io_input_valid),
    .io_iormac(bc_pe_266_io_iormac),
    .io_ve_out(bc_pe_266_io_ve_out),
    .io_ho_out(bc_pe_266_io_ho_out),
    .io_res_out(bc_pe_266_io_res_out)
  );
  bc_pe bc_pe_267 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_267_clock),
    .reset(bc_pe_267_reset),
    .io_ho_input(bc_pe_267_io_ho_input),
    .io_ve_input(bc_pe_267_io_ve_input),
    .io_input_valid(bc_pe_267_io_input_valid),
    .io_iormac(bc_pe_267_io_iormac),
    .io_ve_out(bc_pe_267_io_ve_out),
    .io_ho_out(bc_pe_267_io_ho_out),
    .io_res_out(bc_pe_267_io_res_out)
  );
  bc_pe bc_pe_268 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_268_clock),
    .reset(bc_pe_268_reset),
    .io_ho_input(bc_pe_268_io_ho_input),
    .io_ve_input(bc_pe_268_io_ve_input),
    .io_input_valid(bc_pe_268_io_input_valid),
    .io_iormac(bc_pe_268_io_iormac),
    .io_ve_out(bc_pe_268_io_ve_out),
    .io_ho_out(bc_pe_268_io_ho_out),
    .io_res_out(bc_pe_268_io_res_out)
  );
  bc_pe bc_pe_269 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_269_clock),
    .reset(bc_pe_269_reset),
    .io_ho_input(bc_pe_269_io_ho_input),
    .io_ve_input(bc_pe_269_io_ve_input),
    .io_input_valid(bc_pe_269_io_input_valid),
    .io_iormac(bc_pe_269_io_iormac),
    .io_ve_out(bc_pe_269_io_ve_out),
    .io_ho_out(bc_pe_269_io_ho_out),
    .io_res_out(bc_pe_269_io_res_out)
  );
  bc_pe bc_pe_270 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_270_clock),
    .reset(bc_pe_270_reset),
    .io_ho_input(bc_pe_270_io_ho_input),
    .io_ve_input(bc_pe_270_io_ve_input),
    .io_input_valid(bc_pe_270_io_input_valid),
    .io_iormac(bc_pe_270_io_iormac),
    .io_ve_out(bc_pe_270_io_ve_out),
    .io_ho_out(bc_pe_270_io_ho_out),
    .io_res_out(bc_pe_270_io_res_out)
  );
  bc_pe bc_pe_271 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_271_clock),
    .reset(bc_pe_271_reset),
    .io_ho_input(bc_pe_271_io_ho_input),
    .io_ve_input(bc_pe_271_io_ve_input),
    .io_input_valid(bc_pe_271_io_input_valid),
    .io_iormac(bc_pe_271_io_iormac),
    .io_ve_out(bc_pe_271_io_ve_out),
    .io_ho_out(bc_pe_271_io_ho_out),
    .io_res_out(bc_pe_271_io_res_out)
  );
  bc_pe bc_pe_272 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_272_clock),
    .reset(bc_pe_272_reset),
    .io_ho_input(bc_pe_272_io_ho_input),
    .io_ve_input(bc_pe_272_io_ve_input),
    .io_input_valid(bc_pe_272_io_input_valid),
    .io_iormac(bc_pe_272_io_iormac),
    .io_ve_out(bc_pe_272_io_ve_out),
    .io_ho_out(bc_pe_272_io_ho_out),
    .io_res_out(bc_pe_272_io_res_out)
  );
  bc_pe bc_pe_273 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_273_clock),
    .reset(bc_pe_273_reset),
    .io_ho_input(bc_pe_273_io_ho_input),
    .io_ve_input(bc_pe_273_io_ve_input),
    .io_input_valid(bc_pe_273_io_input_valid),
    .io_iormac(bc_pe_273_io_iormac),
    .io_ve_out(bc_pe_273_io_ve_out),
    .io_ho_out(bc_pe_273_io_ho_out),
    .io_res_out(bc_pe_273_io_res_out)
  );
  bc_pe bc_pe_274 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_274_clock),
    .reset(bc_pe_274_reset),
    .io_ho_input(bc_pe_274_io_ho_input),
    .io_ve_input(bc_pe_274_io_ve_input),
    .io_input_valid(bc_pe_274_io_input_valid),
    .io_iormac(bc_pe_274_io_iormac),
    .io_ve_out(bc_pe_274_io_ve_out),
    .io_ho_out(bc_pe_274_io_ho_out),
    .io_res_out(bc_pe_274_io_res_out)
  );
  bc_pe bc_pe_275 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_275_clock),
    .reset(bc_pe_275_reset),
    .io_ho_input(bc_pe_275_io_ho_input),
    .io_ve_input(bc_pe_275_io_ve_input),
    .io_input_valid(bc_pe_275_io_input_valid),
    .io_iormac(bc_pe_275_io_iormac),
    .io_ve_out(bc_pe_275_io_ve_out),
    .io_ho_out(bc_pe_275_io_ho_out),
    .io_res_out(bc_pe_275_io_res_out)
  );
  bc_pe bc_pe_276 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_276_clock),
    .reset(bc_pe_276_reset),
    .io_ho_input(bc_pe_276_io_ho_input),
    .io_ve_input(bc_pe_276_io_ve_input),
    .io_input_valid(bc_pe_276_io_input_valid),
    .io_iormac(bc_pe_276_io_iormac),
    .io_ve_out(bc_pe_276_io_ve_out),
    .io_ho_out(bc_pe_276_io_ho_out),
    .io_res_out(bc_pe_276_io_res_out)
  );
  bc_pe bc_pe_277 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_277_clock),
    .reset(bc_pe_277_reset),
    .io_ho_input(bc_pe_277_io_ho_input),
    .io_ve_input(bc_pe_277_io_ve_input),
    .io_input_valid(bc_pe_277_io_input_valid),
    .io_iormac(bc_pe_277_io_iormac),
    .io_ve_out(bc_pe_277_io_ve_out),
    .io_ho_out(bc_pe_277_io_ho_out),
    .io_res_out(bc_pe_277_io_res_out)
  );
  bc_pe bc_pe_278 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_278_clock),
    .reset(bc_pe_278_reset),
    .io_ho_input(bc_pe_278_io_ho_input),
    .io_ve_input(bc_pe_278_io_ve_input),
    .io_input_valid(bc_pe_278_io_input_valid),
    .io_iormac(bc_pe_278_io_iormac),
    .io_ve_out(bc_pe_278_io_ve_out),
    .io_ho_out(bc_pe_278_io_ho_out),
    .io_res_out(bc_pe_278_io_res_out)
  );
  bc_pe bc_pe_279 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_279_clock),
    .reset(bc_pe_279_reset),
    .io_ho_input(bc_pe_279_io_ho_input),
    .io_ve_input(bc_pe_279_io_ve_input),
    .io_input_valid(bc_pe_279_io_input_valid),
    .io_iormac(bc_pe_279_io_iormac),
    .io_ve_out(bc_pe_279_io_ve_out),
    .io_ho_out(bc_pe_279_io_ho_out),
    .io_res_out(bc_pe_279_io_res_out)
  );
  bc_pe bc_pe_280 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_280_clock),
    .reset(bc_pe_280_reset),
    .io_ho_input(bc_pe_280_io_ho_input),
    .io_ve_input(bc_pe_280_io_ve_input),
    .io_input_valid(bc_pe_280_io_input_valid),
    .io_iormac(bc_pe_280_io_iormac),
    .io_ve_out(bc_pe_280_io_ve_out),
    .io_ho_out(bc_pe_280_io_ho_out),
    .io_res_out(bc_pe_280_io_res_out)
  );
  bc_pe bc_pe_281 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_281_clock),
    .reset(bc_pe_281_reset),
    .io_ho_input(bc_pe_281_io_ho_input),
    .io_ve_input(bc_pe_281_io_ve_input),
    .io_input_valid(bc_pe_281_io_input_valid),
    .io_iormac(bc_pe_281_io_iormac),
    .io_ve_out(bc_pe_281_io_ve_out),
    .io_ho_out(bc_pe_281_io_ho_out),
    .io_res_out(bc_pe_281_io_res_out)
  );
  bc_pe bc_pe_282 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_282_clock),
    .reset(bc_pe_282_reset),
    .io_ho_input(bc_pe_282_io_ho_input),
    .io_ve_input(bc_pe_282_io_ve_input),
    .io_input_valid(bc_pe_282_io_input_valid),
    .io_iormac(bc_pe_282_io_iormac),
    .io_ve_out(bc_pe_282_io_ve_out),
    .io_ho_out(bc_pe_282_io_ho_out),
    .io_res_out(bc_pe_282_io_res_out)
  );
  bc_pe bc_pe_283 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_283_clock),
    .reset(bc_pe_283_reset),
    .io_ho_input(bc_pe_283_io_ho_input),
    .io_ve_input(bc_pe_283_io_ve_input),
    .io_input_valid(bc_pe_283_io_input_valid),
    .io_iormac(bc_pe_283_io_iormac),
    .io_ve_out(bc_pe_283_io_ve_out),
    .io_ho_out(bc_pe_283_io_ho_out),
    .io_res_out(bc_pe_283_io_res_out)
  );
  bc_pe bc_pe_284 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_284_clock),
    .reset(bc_pe_284_reset),
    .io_ho_input(bc_pe_284_io_ho_input),
    .io_ve_input(bc_pe_284_io_ve_input),
    .io_input_valid(bc_pe_284_io_input_valid),
    .io_iormac(bc_pe_284_io_iormac),
    .io_ve_out(bc_pe_284_io_ve_out),
    .io_ho_out(bc_pe_284_io_ho_out),
    .io_res_out(bc_pe_284_io_res_out)
  );
  bc_pe bc_pe_285 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_285_clock),
    .reset(bc_pe_285_reset),
    .io_ho_input(bc_pe_285_io_ho_input),
    .io_ve_input(bc_pe_285_io_ve_input),
    .io_input_valid(bc_pe_285_io_input_valid),
    .io_iormac(bc_pe_285_io_iormac),
    .io_ve_out(bc_pe_285_io_ve_out),
    .io_ho_out(bc_pe_285_io_ho_out),
    .io_res_out(bc_pe_285_io_res_out)
  );
  bc_pe bc_pe_286 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_286_clock),
    .reset(bc_pe_286_reset),
    .io_ho_input(bc_pe_286_io_ho_input),
    .io_ve_input(bc_pe_286_io_ve_input),
    .io_input_valid(bc_pe_286_io_input_valid),
    .io_iormac(bc_pe_286_io_iormac),
    .io_ve_out(bc_pe_286_io_ve_out),
    .io_ho_out(bc_pe_286_io_ho_out),
    .io_res_out(bc_pe_286_io_res_out)
  );
  bc_pe bc_pe_287 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_287_clock),
    .reset(bc_pe_287_reset),
    .io_ho_input(bc_pe_287_io_ho_input),
    .io_ve_input(bc_pe_287_io_ve_input),
    .io_input_valid(bc_pe_287_io_input_valid),
    .io_iormac(bc_pe_287_io_iormac),
    .io_ve_out(bc_pe_287_io_ve_out),
    .io_ho_out(bc_pe_287_io_ho_out),
    .io_res_out(bc_pe_287_io_res_out)
  );
  bc_pe bc_pe_288 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_288_clock),
    .reset(bc_pe_288_reset),
    .io_ho_input(bc_pe_288_io_ho_input),
    .io_ve_input(bc_pe_288_io_ve_input),
    .io_input_valid(bc_pe_288_io_input_valid),
    .io_iormac(bc_pe_288_io_iormac),
    .io_ve_out(bc_pe_288_io_ve_out),
    .io_ho_out(bc_pe_288_io_ho_out),
    .io_res_out(bc_pe_288_io_res_out)
  );
  bc_pe bc_pe_289 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_289_clock),
    .reset(bc_pe_289_reset),
    .io_ho_input(bc_pe_289_io_ho_input),
    .io_ve_input(bc_pe_289_io_ve_input),
    .io_input_valid(bc_pe_289_io_input_valid),
    .io_iormac(bc_pe_289_io_iormac),
    .io_ve_out(bc_pe_289_io_ve_out),
    .io_ho_out(bc_pe_289_io_ho_out),
    .io_res_out(bc_pe_289_io_res_out)
  );
  bc_pe bc_pe_290 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_290_clock),
    .reset(bc_pe_290_reset),
    .io_ho_input(bc_pe_290_io_ho_input),
    .io_ve_input(bc_pe_290_io_ve_input),
    .io_input_valid(bc_pe_290_io_input_valid),
    .io_iormac(bc_pe_290_io_iormac),
    .io_ve_out(bc_pe_290_io_ve_out),
    .io_ho_out(bc_pe_290_io_ho_out),
    .io_res_out(bc_pe_290_io_res_out)
  );
  bc_pe bc_pe_291 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_291_clock),
    .reset(bc_pe_291_reset),
    .io_ho_input(bc_pe_291_io_ho_input),
    .io_ve_input(bc_pe_291_io_ve_input),
    .io_input_valid(bc_pe_291_io_input_valid),
    .io_iormac(bc_pe_291_io_iormac),
    .io_ve_out(bc_pe_291_io_ve_out),
    .io_ho_out(bc_pe_291_io_ho_out),
    .io_res_out(bc_pe_291_io_res_out)
  );
  bc_pe bc_pe_292 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_292_clock),
    .reset(bc_pe_292_reset),
    .io_ho_input(bc_pe_292_io_ho_input),
    .io_ve_input(bc_pe_292_io_ve_input),
    .io_input_valid(bc_pe_292_io_input_valid),
    .io_iormac(bc_pe_292_io_iormac),
    .io_ve_out(bc_pe_292_io_ve_out),
    .io_ho_out(bc_pe_292_io_ho_out),
    .io_res_out(bc_pe_292_io_res_out)
  );
  bc_pe bc_pe_293 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_293_clock),
    .reset(bc_pe_293_reset),
    .io_ho_input(bc_pe_293_io_ho_input),
    .io_ve_input(bc_pe_293_io_ve_input),
    .io_input_valid(bc_pe_293_io_input_valid),
    .io_iormac(bc_pe_293_io_iormac),
    .io_ve_out(bc_pe_293_io_ve_out),
    .io_ho_out(bc_pe_293_io_ho_out),
    .io_res_out(bc_pe_293_io_res_out)
  );
  bc_pe bc_pe_294 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_294_clock),
    .reset(bc_pe_294_reset),
    .io_ho_input(bc_pe_294_io_ho_input),
    .io_ve_input(bc_pe_294_io_ve_input),
    .io_input_valid(bc_pe_294_io_input_valid),
    .io_iormac(bc_pe_294_io_iormac),
    .io_ve_out(bc_pe_294_io_ve_out),
    .io_ho_out(bc_pe_294_io_ho_out),
    .io_res_out(bc_pe_294_io_res_out)
  );
  bc_pe bc_pe_295 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_295_clock),
    .reset(bc_pe_295_reset),
    .io_ho_input(bc_pe_295_io_ho_input),
    .io_ve_input(bc_pe_295_io_ve_input),
    .io_input_valid(bc_pe_295_io_input_valid),
    .io_iormac(bc_pe_295_io_iormac),
    .io_ve_out(bc_pe_295_io_ve_out),
    .io_ho_out(bc_pe_295_io_ho_out),
    .io_res_out(bc_pe_295_io_res_out)
  );
  bc_pe bc_pe_296 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_296_clock),
    .reset(bc_pe_296_reset),
    .io_ho_input(bc_pe_296_io_ho_input),
    .io_ve_input(bc_pe_296_io_ve_input),
    .io_input_valid(bc_pe_296_io_input_valid),
    .io_iormac(bc_pe_296_io_iormac),
    .io_ve_out(bc_pe_296_io_ve_out),
    .io_ho_out(bc_pe_296_io_ho_out),
    .io_res_out(bc_pe_296_io_res_out)
  );
  bc_pe bc_pe_297 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_297_clock),
    .reset(bc_pe_297_reset),
    .io_ho_input(bc_pe_297_io_ho_input),
    .io_ve_input(bc_pe_297_io_ve_input),
    .io_input_valid(bc_pe_297_io_input_valid),
    .io_iormac(bc_pe_297_io_iormac),
    .io_ve_out(bc_pe_297_io_ve_out),
    .io_ho_out(bc_pe_297_io_ho_out),
    .io_res_out(bc_pe_297_io_res_out)
  );
  bc_pe bc_pe_298 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_298_clock),
    .reset(bc_pe_298_reset),
    .io_ho_input(bc_pe_298_io_ho_input),
    .io_ve_input(bc_pe_298_io_ve_input),
    .io_input_valid(bc_pe_298_io_input_valid),
    .io_iormac(bc_pe_298_io_iormac),
    .io_ve_out(bc_pe_298_io_ve_out),
    .io_ho_out(bc_pe_298_io_ho_out),
    .io_res_out(bc_pe_298_io_res_out)
  );
  bc_pe bc_pe_299 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_299_clock),
    .reset(bc_pe_299_reset),
    .io_ho_input(bc_pe_299_io_ho_input),
    .io_ve_input(bc_pe_299_io_ve_input),
    .io_input_valid(bc_pe_299_io_input_valid),
    .io_iormac(bc_pe_299_io_iormac),
    .io_ve_out(bc_pe_299_io_ve_out),
    .io_ho_out(bc_pe_299_io_ho_out),
    .io_res_out(bc_pe_299_io_res_out)
  );
  bc_pe bc_pe_300 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_300_clock),
    .reset(bc_pe_300_reset),
    .io_ho_input(bc_pe_300_io_ho_input),
    .io_ve_input(bc_pe_300_io_ve_input),
    .io_input_valid(bc_pe_300_io_input_valid),
    .io_iormac(bc_pe_300_io_iormac),
    .io_ve_out(bc_pe_300_io_ve_out),
    .io_ho_out(bc_pe_300_io_ho_out),
    .io_res_out(bc_pe_300_io_res_out)
  );
  bc_pe bc_pe_301 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_301_clock),
    .reset(bc_pe_301_reset),
    .io_ho_input(bc_pe_301_io_ho_input),
    .io_ve_input(bc_pe_301_io_ve_input),
    .io_input_valid(bc_pe_301_io_input_valid),
    .io_iormac(bc_pe_301_io_iormac),
    .io_ve_out(bc_pe_301_io_ve_out),
    .io_ho_out(bc_pe_301_io_ho_out),
    .io_res_out(bc_pe_301_io_res_out)
  );
  bc_pe bc_pe_302 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_302_clock),
    .reset(bc_pe_302_reset),
    .io_ho_input(bc_pe_302_io_ho_input),
    .io_ve_input(bc_pe_302_io_ve_input),
    .io_input_valid(bc_pe_302_io_input_valid),
    .io_iormac(bc_pe_302_io_iormac),
    .io_ve_out(bc_pe_302_io_ve_out),
    .io_ho_out(bc_pe_302_io_ho_out),
    .io_res_out(bc_pe_302_io_res_out)
  );
  bc_pe bc_pe_303 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_303_clock),
    .reset(bc_pe_303_reset),
    .io_ho_input(bc_pe_303_io_ho_input),
    .io_ve_input(bc_pe_303_io_ve_input),
    .io_input_valid(bc_pe_303_io_input_valid),
    .io_iormac(bc_pe_303_io_iormac),
    .io_ve_out(bc_pe_303_io_ve_out),
    .io_ho_out(bc_pe_303_io_ho_out),
    .io_res_out(bc_pe_303_io_res_out)
  );
  bc_pe bc_pe_304 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_304_clock),
    .reset(bc_pe_304_reset),
    .io_ho_input(bc_pe_304_io_ho_input),
    .io_ve_input(bc_pe_304_io_ve_input),
    .io_input_valid(bc_pe_304_io_input_valid),
    .io_iormac(bc_pe_304_io_iormac),
    .io_ve_out(bc_pe_304_io_ve_out),
    .io_ho_out(bc_pe_304_io_ho_out),
    .io_res_out(bc_pe_304_io_res_out)
  );
  bc_pe bc_pe_305 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_305_clock),
    .reset(bc_pe_305_reset),
    .io_ho_input(bc_pe_305_io_ho_input),
    .io_ve_input(bc_pe_305_io_ve_input),
    .io_input_valid(bc_pe_305_io_input_valid),
    .io_iormac(bc_pe_305_io_iormac),
    .io_ve_out(bc_pe_305_io_ve_out),
    .io_ho_out(bc_pe_305_io_ho_out),
    .io_res_out(bc_pe_305_io_res_out)
  );
  bc_pe bc_pe_306 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_306_clock),
    .reset(bc_pe_306_reset),
    .io_ho_input(bc_pe_306_io_ho_input),
    .io_ve_input(bc_pe_306_io_ve_input),
    .io_input_valid(bc_pe_306_io_input_valid),
    .io_iormac(bc_pe_306_io_iormac),
    .io_ve_out(bc_pe_306_io_ve_out),
    .io_ho_out(bc_pe_306_io_ho_out),
    .io_res_out(bc_pe_306_io_res_out)
  );
  bc_pe bc_pe_307 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_307_clock),
    .reset(bc_pe_307_reset),
    .io_ho_input(bc_pe_307_io_ho_input),
    .io_ve_input(bc_pe_307_io_ve_input),
    .io_input_valid(bc_pe_307_io_input_valid),
    .io_iormac(bc_pe_307_io_iormac),
    .io_ve_out(bc_pe_307_io_ve_out),
    .io_ho_out(bc_pe_307_io_ho_out),
    .io_res_out(bc_pe_307_io_res_out)
  );
  bc_pe bc_pe_308 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_308_clock),
    .reset(bc_pe_308_reset),
    .io_ho_input(bc_pe_308_io_ho_input),
    .io_ve_input(bc_pe_308_io_ve_input),
    .io_input_valid(bc_pe_308_io_input_valid),
    .io_iormac(bc_pe_308_io_iormac),
    .io_ve_out(bc_pe_308_io_ve_out),
    .io_ho_out(bc_pe_308_io_ho_out),
    .io_res_out(bc_pe_308_io_res_out)
  );
  bc_pe bc_pe_309 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_309_clock),
    .reset(bc_pe_309_reset),
    .io_ho_input(bc_pe_309_io_ho_input),
    .io_ve_input(bc_pe_309_io_ve_input),
    .io_input_valid(bc_pe_309_io_input_valid),
    .io_iormac(bc_pe_309_io_iormac),
    .io_ve_out(bc_pe_309_io_ve_out),
    .io_ho_out(bc_pe_309_io_ho_out),
    .io_res_out(bc_pe_309_io_res_out)
  );
  bc_pe bc_pe_310 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_310_clock),
    .reset(bc_pe_310_reset),
    .io_ho_input(bc_pe_310_io_ho_input),
    .io_ve_input(bc_pe_310_io_ve_input),
    .io_input_valid(bc_pe_310_io_input_valid),
    .io_iormac(bc_pe_310_io_iormac),
    .io_ve_out(bc_pe_310_io_ve_out),
    .io_ho_out(bc_pe_310_io_ho_out),
    .io_res_out(bc_pe_310_io_res_out)
  );
  bc_pe bc_pe_311 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_311_clock),
    .reset(bc_pe_311_reset),
    .io_ho_input(bc_pe_311_io_ho_input),
    .io_ve_input(bc_pe_311_io_ve_input),
    .io_input_valid(bc_pe_311_io_input_valid),
    .io_iormac(bc_pe_311_io_iormac),
    .io_ve_out(bc_pe_311_io_ve_out),
    .io_ho_out(bc_pe_311_io_ho_out),
    .io_res_out(bc_pe_311_io_res_out)
  );
  bc_pe bc_pe_312 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_312_clock),
    .reset(bc_pe_312_reset),
    .io_ho_input(bc_pe_312_io_ho_input),
    .io_ve_input(bc_pe_312_io_ve_input),
    .io_input_valid(bc_pe_312_io_input_valid),
    .io_iormac(bc_pe_312_io_iormac),
    .io_ve_out(bc_pe_312_io_ve_out),
    .io_ho_out(bc_pe_312_io_ho_out),
    .io_res_out(bc_pe_312_io_res_out)
  );
  bc_pe bc_pe_313 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_313_clock),
    .reset(bc_pe_313_reset),
    .io_ho_input(bc_pe_313_io_ho_input),
    .io_ve_input(bc_pe_313_io_ve_input),
    .io_input_valid(bc_pe_313_io_input_valid),
    .io_iormac(bc_pe_313_io_iormac),
    .io_ve_out(bc_pe_313_io_ve_out),
    .io_ho_out(bc_pe_313_io_ho_out),
    .io_res_out(bc_pe_313_io_res_out)
  );
  bc_pe bc_pe_314 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_314_clock),
    .reset(bc_pe_314_reset),
    .io_ho_input(bc_pe_314_io_ho_input),
    .io_ve_input(bc_pe_314_io_ve_input),
    .io_input_valid(bc_pe_314_io_input_valid),
    .io_iormac(bc_pe_314_io_iormac),
    .io_ve_out(bc_pe_314_io_ve_out),
    .io_ho_out(bc_pe_314_io_ho_out),
    .io_res_out(bc_pe_314_io_res_out)
  );
  bc_pe bc_pe_315 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_315_clock),
    .reset(bc_pe_315_reset),
    .io_ho_input(bc_pe_315_io_ho_input),
    .io_ve_input(bc_pe_315_io_ve_input),
    .io_input_valid(bc_pe_315_io_input_valid),
    .io_iormac(bc_pe_315_io_iormac),
    .io_ve_out(bc_pe_315_io_ve_out),
    .io_ho_out(bc_pe_315_io_ho_out),
    .io_res_out(bc_pe_315_io_res_out)
  );
  bc_pe bc_pe_316 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_316_clock),
    .reset(bc_pe_316_reset),
    .io_ho_input(bc_pe_316_io_ho_input),
    .io_ve_input(bc_pe_316_io_ve_input),
    .io_input_valid(bc_pe_316_io_input_valid),
    .io_iormac(bc_pe_316_io_iormac),
    .io_ve_out(bc_pe_316_io_ve_out),
    .io_ho_out(bc_pe_316_io_ho_out),
    .io_res_out(bc_pe_316_io_res_out)
  );
  bc_pe bc_pe_317 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_317_clock),
    .reset(bc_pe_317_reset),
    .io_ho_input(bc_pe_317_io_ho_input),
    .io_ve_input(bc_pe_317_io_ve_input),
    .io_input_valid(bc_pe_317_io_input_valid),
    .io_iormac(bc_pe_317_io_iormac),
    .io_ve_out(bc_pe_317_io_ve_out),
    .io_ho_out(bc_pe_317_io_ho_out),
    .io_res_out(bc_pe_317_io_res_out)
  );
  bc_pe bc_pe_318 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_318_clock),
    .reset(bc_pe_318_reset),
    .io_ho_input(bc_pe_318_io_ho_input),
    .io_ve_input(bc_pe_318_io_ve_input),
    .io_input_valid(bc_pe_318_io_input_valid),
    .io_iormac(bc_pe_318_io_iormac),
    .io_ve_out(bc_pe_318_io_ve_out),
    .io_ho_out(bc_pe_318_io_ho_out),
    .io_res_out(bc_pe_318_io_res_out)
  );
  bc_pe bc_pe_319 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_319_clock),
    .reset(bc_pe_319_reset),
    .io_ho_input(bc_pe_319_io_ho_input),
    .io_ve_input(bc_pe_319_io_ve_input),
    .io_input_valid(bc_pe_319_io_input_valid),
    .io_iormac(bc_pe_319_io_iormac),
    .io_ve_out(bc_pe_319_io_ve_out),
    .io_ho_out(bc_pe_319_io_ho_out),
    .io_res_out(bc_pe_319_io_res_out)
  );
  bc_pe bc_pe_320 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_320_clock),
    .reset(bc_pe_320_reset),
    .io_ho_input(bc_pe_320_io_ho_input),
    .io_ve_input(bc_pe_320_io_ve_input),
    .io_input_valid(bc_pe_320_io_input_valid),
    .io_iormac(bc_pe_320_io_iormac),
    .io_ve_out(bc_pe_320_io_ve_out),
    .io_ho_out(bc_pe_320_io_ho_out),
    .io_res_out(bc_pe_320_io_res_out)
  );
  bc_pe bc_pe_321 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_321_clock),
    .reset(bc_pe_321_reset),
    .io_ho_input(bc_pe_321_io_ho_input),
    .io_ve_input(bc_pe_321_io_ve_input),
    .io_input_valid(bc_pe_321_io_input_valid),
    .io_iormac(bc_pe_321_io_iormac),
    .io_ve_out(bc_pe_321_io_ve_out),
    .io_ho_out(bc_pe_321_io_ho_out),
    .io_res_out(bc_pe_321_io_res_out)
  );
  bc_pe bc_pe_322 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_322_clock),
    .reset(bc_pe_322_reset),
    .io_ho_input(bc_pe_322_io_ho_input),
    .io_ve_input(bc_pe_322_io_ve_input),
    .io_input_valid(bc_pe_322_io_input_valid),
    .io_iormac(bc_pe_322_io_iormac),
    .io_ve_out(bc_pe_322_io_ve_out),
    .io_ho_out(bc_pe_322_io_ho_out),
    .io_res_out(bc_pe_322_io_res_out)
  );
  bc_pe bc_pe_323 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_323_clock),
    .reset(bc_pe_323_reset),
    .io_ho_input(bc_pe_323_io_ho_input),
    .io_ve_input(bc_pe_323_io_ve_input),
    .io_input_valid(bc_pe_323_io_input_valid),
    .io_iormac(bc_pe_323_io_iormac),
    .io_ve_out(bc_pe_323_io_ve_out),
    .io_ho_out(bc_pe_323_io_ho_out),
    .io_res_out(bc_pe_323_io_res_out)
  );
  bc_pe bc_pe_324 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_324_clock),
    .reset(bc_pe_324_reset),
    .io_ho_input(bc_pe_324_io_ho_input),
    .io_ve_input(bc_pe_324_io_ve_input),
    .io_input_valid(bc_pe_324_io_input_valid),
    .io_iormac(bc_pe_324_io_iormac),
    .io_ve_out(bc_pe_324_io_ve_out),
    .io_ho_out(bc_pe_324_io_ho_out),
    .io_res_out(bc_pe_324_io_res_out)
  );
  bc_pe bc_pe_325 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_325_clock),
    .reset(bc_pe_325_reset),
    .io_ho_input(bc_pe_325_io_ho_input),
    .io_ve_input(bc_pe_325_io_ve_input),
    .io_input_valid(bc_pe_325_io_input_valid),
    .io_iormac(bc_pe_325_io_iormac),
    .io_ve_out(bc_pe_325_io_ve_out),
    .io_ho_out(bc_pe_325_io_ho_out),
    .io_res_out(bc_pe_325_io_res_out)
  );
  bc_pe bc_pe_326 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_326_clock),
    .reset(bc_pe_326_reset),
    .io_ho_input(bc_pe_326_io_ho_input),
    .io_ve_input(bc_pe_326_io_ve_input),
    .io_input_valid(bc_pe_326_io_input_valid),
    .io_iormac(bc_pe_326_io_iormac),
    .io_ve_out(bc_pe_326_io_ve_out),
    .io_ho_out(bc_pe_326_io_ho_out),
    .io_res_out(bc_pe_326_io_res_out)
  );
  bc_pe bc_pe_327 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_327_clock),
    .reset(bc_pe_327_reset),
    .io_ho_input(bc_pe_327_io_ho_input),
    .io_ve_input(bc_pe_327_io_ve_input),
    .io_input_valid(bc_pe_327_io_input_valid),
    .io_iormac(bc_pe_327_io_iormac),
    .io_ve_out(bc_pe_327_io_ve_out),
    .io_ho_out(bc_pe_327_io_ho_out),
    .io_res_out(bc_pe_327_io_res_out)
  );
  bc_pe bc_pe_328 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_328_clock),
    .reset(bc_pe_328_reset),
    .io_ho_input(bc_pe_328_io_ho_input),
    .io_ve_input(bc_pe_328_io_ve_input),
    .io_input_valid(bc_pe_328_io_input_valid),
    .io_iormac(bc_pe_328_io_iormac),
    .io_ve_out(bc_pe_328_io_ve_out),
    .io_ho_out(bc_pe_328_io_ho_out),
    .io_res_out(bc_pe_328_io_res_out)
  );
  bc_pe bc_pe_329 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_329_clock),
    .reset(bc_pe_329_reset),
    .io_ho_input(bc_pe_329_io_ho_input),
    .io_ve_input(bc_pe_329_io_ve_input),
    .io_input_valid(bc_pe_329_io_input_valid),
    .io_iormac(bc_pe_329_io_iormac),
    .io_ve_out(bc_pe_329_io_ve_out),
    .io_ho_out(bc_pe_329_io_ho_out),
    .io_res_out(bc_pe_329_io_res_out)
  );
  bc_pe bc_pe_330 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_330_clock),
    .reset(bc_pe_330_reset),
    .io_ho_input(bc_pe_330_io_ho_input),
    .io_ve_input(bc_pe_330_io_ve_input),
    .io_input_valid(bc_pe_330_io_input_valid),
    .io_iormac(bc_pe_330_io_iormac),
    .io_ve_out(bc_pe_330_io_ve_out),
    .io_ho_out(bc_pe_330_io_ho_out),
    .io_res_out(bc_pe_330_io_res_out)
  );
  bc_pe bc_pe_331 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_331_clock),
    .reset(bc_pe_331_reset),
    .io_ho_input(bc_pe_331_io_ho_input),
    .io_ve_input(bc_pe_331_io_ve_input),
    .io_input_valid(bc_pe_331_io_input_valid),
    .io_iormac(bc_pe_331_io_iormac),
    .io_ve_out(bc_pe_331_io_ve_out),
    .io_ho_out(bc_pe_331_io_ho_out),
    .io_res_out(bc_pe_331_io_res_out)
  );
  bc_pe bc_pe_332 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_332_clock),
    .reset(bc_pe_332_reset),
    .io_ho_input(bc_pe_332_io_ho_input),
    .io_ve_input(bc_pe_332_io_ve_input),
    .io_input_valid(bc_pe_332_io_input_valid),
    .io_iormac(bc_pe_332_io_iormac),
    .io_ve_out(bc_pe_332_io_ve_out),
    .io_ho_out(bc_pe_332_io_ho_out),
    .io_res_out(bc_pe_332_io_res_out)
  );
  bc_pe bc_pe_333 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_333_clock),
    .reset(bc_pe_333_reset),
    .io_ho_input(bc_pe_333_io_ho_input),
    .io_ve_input(bc_pe_333_io_ve_input),
    .io_input_valid(bc_pe_333_io_input_valid),
    .io_iormac(bc_pe_333_io_iormac),
    .io_ve_out(bc_pe_333_io_ve_out),
    .io_ho_out(bc_pe_333_io_ho_out),
    .io_res_out(bc_pe_333_io_res_out)
  );
  bc_pe bc_pe_334 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_334_clock),
    .reset(bc_pe_334_reset),
    .io_ho_input(bc_pe_334_io_ho_input),
    .io_ve_input(bc_pe_334_io_ve_input),
    .io_input_valid(bc_pe_334_io_input_valid),
    .io_iormac(bc_pe_334_io_iormac),
    .io_ve_out(bc_pe_334_io_ve_out),
    .io_ho_out(bc_pe_334_io_ho_out),
    .io_res_out(bc_pe_334_io_res_out)
  );
  bc_pe bc_pe_335 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_335_clock),
    .reset(bc_pe_335_reset),
    .io_ho_input(bc_pe_335_io_ho_input),
    .io_ve_input(bc_pe_335_io_ve_input),
    .io_input_valid(bc_pe_335_io_input_valid),
    .io_iormac(bc_pe_335_io_iormac),
    .io_ve_out(bc_pe_335_io_ve_out),
    .io_ho_out(bc_pe_335_io_ho_out),
    .io_res_out(bc_pe_335_io_res_out)
  );
  bc_pe bc_pe_336 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_336_clock),
    .reset(bc_pe_336_reset),
    .io_ho_input(bc_pe_336_io_ho_input),
    .io_ve_input(bc_pe_336_io_ve_input),
    .io_input_valid(bc_pe_336_io_input_valid),
    .io_iormac(bc_pe_336_io_iormac),
    .io_ve_out(bc_pe_336_io_ve_out),
    .io_ho_out(bc_pe_336_io_ho_out),
    .io_res_out(bc_pe_336_io_res_out)
  );
  bc_pe bc_pe_337 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_337_clock),
    .reset(bc_pe_337_reset),
    .io_ho_input(bc_pe_337_io_ho_input),
    .io_ve_input(bc_pe_337_io_ve_input),
    .io_input_valid(bc_pe_337_io_input_valid),
    .io_iormac(bc_pe_337_io_iormac),
    .io_ve_out(bc_pe_337_io_ve_out),
    .io_ho_out(bc_pe_337_io_ho_out),
    .io_res_out(bc_pe_337_io_res_out)
  );
  bc_pe bc_pe_338 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_338_clock),
    .reset(bc_pe_338_reset),
    .io_ho_input(bc_pe_338_io_ho_input),
    .io_ve_input(bc_pe_338_io_ve_input),
    .io_input_valid(bc_pe_338_io_input_valid),
    .io_iormac(bc_pe_338_io_iormac),
    .io_ve_out(bc_pe_338_io_ve_out),
    .io_ho_out(bc_pe_338_io_ho_out),
    .io_res_out(bc_pe_338_io_res_out)
  );
  bc_pe bc_pe_339 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_339_clock),
    .reset(bc_pe_339_reset),
    .io_ho_input(bc_pe_339_io_ho_input),
    .io_ve_input(bc_pe_339_io_ve_input),
    .io_input_valid(bc_pe_339_io_input_valid),
    .io_iormac(bc_pe_339_io_iormac),
    .io_ve_out(bc_pe_339_io_ve_out),
    .io_ho_out(bc_pe_339_io_ho_out),
    .io_res_out(bc_pe_339_io_res_out)
  );
  bc_pe bc_pe_340 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_340_clock),
    .reset(bc_pe_340_reset),
    .io_ho_input(bc_pe_340_io_ho_input),
    .io_ve_input(bc_pe_340_io_ve_input),
    .io_input_valid(bc_pe_340_io_input_valid),
    .io_iormac(bc_pe_340_io_iormac),
    .io_ve_out(bc_pe_340_io_ve_out),
    .io_ho_out(bc_pe_340_io_ho_out),
    .io_res_out(bc_pe_340_io_res_out)
  );
  bc_pe bc_pe_341 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_341_clock),
    .reset(bc_pe_341_reset),
    .io_ho_input(bc_pe_341_io_ho_input),
    .io_ve_input(bc_pe_341_io_ve_input),
    .io_input_valid(bc_pe_341_io_input_valid),
    .io_iormac(bc_pe_341_io_iormac),
    .io_ve_out(bc_pe_341_io_ve_out),
    .io_ho_out(bc_pe_341_io_ho_out),
    .io_res_out(bc_pe_341_io_res_out)
  );
  bc_pe bc_pe_342 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_342_clock),
    .reset(bc_pe_342_reset),
    .io_ho_input(bc_pe_342_io_ho_input),
    .io_ve_input(bc_pe_342_io_ve_input),
    .io_input_valid(bc_pe_342_io_input_valid),
    .io_iormac(bc_pe_342_io_iormac),
    .io_ve_out(bc_pe_342_io_ve_out),
    .io_ho_out(bc_pe_342_io_ho_out),
    .io_res_out(bc_pe_342_io_res_out)
  );
  bc_pe bc_pe_343 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_343_clock),
    .reset(bc_pe_343_reset),
    .io_ho_input(bc_pe_343_io_ho_input),
    .io_ve_input(bc_pe_343_io_ve_input),
    .io_input_valid(bc_pe_343_io_input_valid),
    .io_iormac(bc_pe_343_io_iormac),
    .io_ve_out(bc_pe_343_io_ve_out),
    .io_ho_out(bc_pe_343_io_ho_out),
    .io_res_out(bc_pe_343_io_res_out)
  );
  bc_pe bc_pe_344 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_344_clock),
    .reset(bc_pe_344_reset),
    .io_ho_input(bc_pe_344_io_ho_input),
    .io_ve_input(bc_pe_344_io_ve_input),
    .io_input_valid(bc_pe_344_io_input_valid),
    .io_iormac(bc_pe_344_io_iormac),
    .io_ve_out(bc_pe_344_io_ve_out),
    .io_ho_out(bc_pe_344_io_ho_out),
    .io_res_out(bc_pe_344_io_res_out)
  );
  bc_pe bc_pe_345 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_345_clock),
    .reset(bc_pe_345_reset),
    .io_ho_input(bc_pe_345_io_ho_input),
    .io_ve_input(bc_pe_345_io_ve_input),
    .io_input_valid(bc_pe_345_io_input_valid),
    .io_iormac(bc_pe_345_io_iormac),
    .io_ve_out(bc_pe_345_io_ve_out),
    .io_ho_out(bc_pe_345_io_ho_out),
    .io_res_out(bc_pe_345_io_res_out)
  );
  bc_pe bc_pe_346 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_346_clock),
    .reset(bc_pe_346_reset),
    .io_ho_input(bc_pe_346_io_ho_input),
    .io_ve_input(bc_pe_346_io_ve_input),
    .io_input_valid(bc_pe_346_io_input_valid),
    .io_iormac(bc_pe_346_io_iormac),
    .io_ve_out(bc_pe_346_io_ve_out),
    .io_ho_out(bc_pe_346_io_ho_out),
    .io_res_out(bc_pe_346_io_res_out)
  );
  bc_pe bc_pe_347 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_347_clock),
    .reset(bc_pe_347_reset),
    .io_ho_input(bc_pe_347_io_ho_input),
    .io_ve_input(bc_pe_347_io_ve_input),
    .io_input_valid(bc_pe_347_io_input_valid),
    .io_iormac(bc_pe_347_io_iormac),
    .io_ve_out(bc_pe_347_io_ve_out),
    .io_ho_out(bc_pe_347_io_ho_out),
    .io_res_out(bc_pe_347_io_res_out)
  );
  bc_pe bc_pe_348 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_348_clock),
    .reset(bc_pe_348_reset),
    .io_ho_input(bc_pe_348_io_ho_input),
    .io_ve_input(bc_pe_348_io_ve_input),
    .io_input_valid(bc_pe_348_io_input_valid),
    .io_iormac(bc_pe_348_io_iormac),
    .io_ve_out(bc_pe_348_io_ve_out),
    .io_ho_out(bc_pe_348_io_ho_out),
    .io_res_out(bc_pe_348_io_res_out)
  );
  bc_pe bc_pe_349 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_349_clock),
    .reset(bc_pe_349_reset),
    .io_ho_input(bc_pe_349_io_ho_input),
    .io_ve_input(bc_pe_349_io_ve_input),
    .io_input_valid(bc_pe_349_io_input_valid),
    .io_iormac(bc_pe_349_io_iormac),
    .io_ve_out(bc_pe_349_io_ve_out),
    .io_ho_out(bc_pe_349_io_ho_out),
    .io_res_out(bc_pe_349_io_res_out)
  );
  bc_pe bc_pe_350 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_350_clock),
    .reset(bc_pe_350_reset),
    .io_ho_input(bc_pe_350_io_ho_input),
    .io_ve_input(bc_pe_350_io_ve_input),
    .io_input_valid(bc_pe_350_io_input_valid),
    .io_iormac(bc_pe_350_io_iormac),
    .io_ve_out(bc_pe_350_io_ve_out),
    .io_ho_out(bc_pe_350_io_ho_out),
    .io_res_out(bc_pe_350_io_res_out)
  );
  bc_pe bc_pe_351 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_351_clock),
    .reset(bc_pe_351_reset),
    .io_ho_input(bc_pe_351_io_ho_input),
    .io_ve_input(bc_pe_351_io_ve_input),
    .io_input_valid(bc_pe_351_io_input_valid),
    .io_iormac(bc_pe_351_io_iormac),
    .io_ve_out(bc_pe_351_io_ve_out),
    .io_ho_out(bc_pe_351_io_ho_out),
    .io_res_out(bc_pe_351_io_res_out)
  );
  bc_pe bc_pe_352 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_352_clock),
    .reset(bc_pe_352_reset),
    .io_ho_input(bc_pe_352_io_ho_input),
    .io_ve_input(bc_pe_352_io_ve_input),
    .io_input_valid(bc_pe_352_io_input_valid),
    .io_iormac(bc_pe_352_io_iormac),
    .io_ve_out(bc_pe_352_io_ve_out),
    .io_ho_out(bc_pe_352_io_ho_out),
    .io_res_out(bc_pe_352_io_res_out)
  );
  bc_pe bc_pe_353 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_353_clock),
    .reset(bc_pe_353_reset),
    .io_ho_input(bc_pe_353_io_ho_input),
    .io_ve_input(bc_pe_353_io_ve_input),
    .io_input_valid(bc_pe_353_io_input_valid),
    .io_iormac(bc_pe_353_io_iormac),
    .io_ve_out(bc_pe_353_io_ve_out),
    .io_ho_out(bc_pe_353_io_ho_out),
    .io_res_out(bc_pe_353_io_res_out)
  );
  bc_pe bc_pe_354 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_354_clock),
    .reset(bc_pe_354_reset),
    .io_ho_input(bc_pe_354_io_ho_input),
    .io_ve_input(bc_pe_354_io_ve_input),
    .io_input_valid(bc_pe_354_io_input_valid),
    .io_iormac(bc_pe_354_io_iormac),
    .io_ve_out(bc_pe_354_io_ve_out),
    .io_ho_out(bc_pe_354_io_ho_out),
    .io_res_out(bc_pe_354_io_res_out)
  );
  bc_pe bc_pe_355 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_355_clock),
    .reset(bc_pe_355_reset),
    .io_ho_input(bc_pe_355_io_ho_input),
    .io_ve_input(bc_pe_355_io_ve_input),
    .io_input_valid(bc_pe_355_io_input_valid),
    .io_iormac(bc_pe_355_io_iormac),
    .io_ve_out(bc_pe_355_io_ve_out),
    .io_ho_out(bc_pe_355_io_ho_out),
    .io_res_out(bc_pe_355_io_res_out)
  );
  bc_pe bc_pe_356 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_356_clock),
    .reset(bc_pe_356_reset),
    .io_ho_input(bc_pe_356_io_ho_input),
    .io_ve_input(bc_pe_356_io_ve_input),
    .io_input_valid(bc_pe_356_io_input_valid),
    .io_iormac(bc_pe_356_io_iormac),
    .io_ve_out(bc_pe_356_io_ve_out),
    .io_ho_out(bc_pe_356_io_ho_out),
    .io_res_out(bc_pe_356_io_res_out)
  );
  bc_pe bc_pe_357 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_357_clock),
    .reset(bc_pe_357_reset),
    .io_ho_input(bc_pe_357_io_ho_input),
    .io_ve_input(bc_pe_357_io_ve_input),
    .io_input_valid(bc_pe_357_io_input_valid),
    .io_iormac(bc_pe_357_io_iormac),
    .io_ve_out(bc_pe_357_io_ve_out),
    .io_ho_out(bc_pe_357_io_ho_out),
    .io_res_out(bc_pe_357_io_res_out)
  );
  bc_pe bc_pe_358 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_358_clock),
    .reset(bc_pe_358_reset),
    .io_ho_input(bc_pe_358_io_ho_input),
    .io_ve_input(bc_pe_358_io_ve_input),
    .io_input_valid(bc_pe_358_io_input_valid),
    .io_iormac(bc_pe_358_io_iormac),
    .io_ve_out(bc_pe_358_io_ve_out),
    .io_ho_out(bc_pe_358_io_ho_out),
    .io_res_out(bc_pe_358_io_res_out)
  );
  bc_pe bc_pe_359 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_359_clock),
    .reset(bc_pe_359_reset),
    .io_ho_input(bc_pe_359_io_ho_input),
    .io_ve_input(bc_pe_359_io_ve_input),
    .io_input_valid(bc_pe_359_io_input_valid),
    .io_iormac(bc_pe_359_io_iormac),
    .io_ve_out(bc_pe_359_io_ve_out),
    .io_ho_out(bc_pe_359_io_ho_out),
    .io_res_out(bc_pe_359_io_res_out)
  );
  bc_pe bc_pe_360 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_360_clock),
    .reset(bc_pe_360_reset),
    .io_ho_input(bc_pe_360_io_ho_input),
    .io_ve_input(bc_pe_360_io_ve_input),
    .io_input_valid(bc_pe_360_io_input_valid),
    .io_iormac(bc_pe_360_io_iormac),
    .io_ve_out(bc_pe_360_io_ve_out),
    .io_ho_out(bc_pe_360_io_ho_out),
    .io_res_out(bc_pe_360_io_res_out)
  );
  bc_pe bc_pe_361 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_361_clock),
    .reset(bc_pe_361_reset),
    .io_ho_input(bc_pe_361_io_ho_input),
    .io_ve_input(bc_pe_361_io_ve_input),
    .io_input_valid(bc_pe_361_io_input_valid),
    .io_iormac(bc_pe_361_io_iormac),
    .io_ve_out(bc_pe_361_io_ve_out),
    .io_ho_out(bc_pe_361_io_ho_out),
    .io_res_out(bc_pe_361_io_res_out)
  );
  bc_pe bc_pe_362 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_362_clock),
    .reset(bc_pe_362_reset),
    .io_ho_input(bc_pe_362_io_ho_input),
    .io_ve_input(bc_pe_362_io_ve_input),
    .io_input_valid(bc_pe_362_io_input_valid),
    .io_iormac(bc_pe_362_io_iormac),
    .io_ve_out(bc_pe_362_io_ve_out),
    .io_ho_out(bc_pe_362_io_ho_out),
    .io_res_out(bc_pe_362_io_res_out)
  );
  bc_pe bc_pe_363 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_363_clock),
    .reset(bc_pe_363_reset),
    .io_ho_input(bc_pe_363_io_ho_input),
    .io_ve_input(bc_pe_363_io_ve_input),
    .io_input_valid(bc_pe_363_io_input_valid),
    .io_iormac(bc_pe_363_io_iormac),
    .io_ve_out(bc_pe_363_io_ve_out),
    .io_ho_out(bc_pe_363_io_ho_out),
    .io_res_out(bc_pe_363_io_res_out)
  );
  bc_pe bc_pe_364 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_364_clock),
    .reset(bc_pe_364_reset),
    .io_ho_input(bc_pe_364_io_ho_input),
    .io_ve_input(bc_pe_364_io_ve_input),
    .io_input_valid(bc_pe_364_io_input_valid),
    .io_iormac(bc_pe_364_io_iormac),
    .io_ve_out(bc_pe_364_io_ve_out),
    .io_ho_out(bc_pe_364_io_ho_out),
    .io_res_out(bc_pe_364_io_res_out)
  );
  bc_pe bc_pe_365 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_365_clock),
    .reset(bc_pe_365_reset),
    .io_ho_input(bc_pe_365_io_ho_input),
    .io_ve_input(bc_pe_365_io_ve_input),
    .io_input_valid(bc_pe_365_io_input_valid),
    .io_iormac(bc_pe_365_io_iormac),
    .io_ve_out(bc_pe_365_io_ve_out),
    .io_ho_out(bc_pe_365_io_ho_out),
    .io_res_out(bc_pe_365_io_res_out)
  );
  bc_pe bc_pe_366 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_366_clock),
    .reset(bc_pe_366_reset),
    .io_ho_input(bc_pe_366_io_ho_input),
    .io_ve_input(bc_pe_366_io_ve_input),
    .io_input_valid(bc_pe_366_io_input_valid),
    .io_iormac(bc_pe_366_io_iormac),
    .io_ve_out(bc_pe_366_io_ve_out),
    .io_ho_out(bc_pe_366_io_ho_out),
    .io_res_out(bc_pe_366_io_res_out)
  );
  bc_pe bc_pe_367 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_367_clock),
    .reset(bc_pe_367_reset),
    .io_ho_input(bc_pe_367_io_ho_input),
    .io_ve_input(bc_pe_367_io_ve_input),
    .io_input_valid(bc_pe_367_io_input_valid),
    .io_iormac(bc_pe_367_io_iormac),
    .io_ve_out(bc_pe_367_io_ve_out),
    .io_ho_out(bc_pe_367_io_ho_out),
    .io_res_out(bc_pe_367_io_res_out)
  );
  bc_pe bc_pe_368 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_368_clock),
    .reset(bc_pe_368_reset),
    .io_ho_input(bc_pe_368_io_ho_input),
    .io_ve_input(bc_pe_368_io_ve_input),
    .io_input_valid(bc_pe_368_io_input_valid),
    .io_iormac(bc_pe_368_io_iormac),
    .io_ve_out(bc_pe_368_io_ve_out),
    .io_ho_out(bc_pe_368_io_ho_out),
    .io_res_out(bc_pe_368_io_res_out)
  );
  bc_pe bc_pe_369 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_369_clock),
    .reset(bc_pe_369_reset),
    .io_ho_input(bc_pe_369_io_ho_input),
    .io_ve_input(bc_pe_369_io_ve_input),
    .io_input_valid(bc_pe_369_io_input_valid),
    .io_iormac(bc_pe_369_io_iormac),
    .io_ve_out(bc_pe_369_io_ve_out),
    .io_ho_out(bc_pe_369_io_ho_out),
    .io_res_out(bc_pe_369_io_res_out)
  );
  bc_pe bc_pe_370 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_370_clock),
    .reset(bc_pe_370_reset),
    .io_ho_input(bc_pe_370_io_ho_input),
    .io_ve_input(bc_pe_370_io_ve_input),
    .io_input_valid(bc_pe_370_io_input_valid),
    .io_iormac(bc_pe_370_io_iormac),
    .io_ve_out(bc_pe_370_io_ve_out),
    .io_ho_out(bc_pe_370_io_ho_out),
    .io_res_out(bc_pe_370_io_res_out)
  );
  bc_pe bc_pe_371 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_371_clock),
    .reset(bc_pe_371_reset),
    .io_ho_input(bc_pe_371_io_ho_input),
    .io_ve_input(bc_pe_371_io_ve_input),
    .io_input_valid(bc_pe_371_io_input_valid),
    .io_iormac(bc_pe_371_io_iormac),
    .io_ve_out(bc_pe_371_io_ve_out),
    .io_ho_out(bc_pe_371_io_ho_out),
    .io_res_out(bc_pe_371_io_res_out)
  );
  bc_pe bc_pe_372 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_372_clock),
    .reset(bc_pe_372_reset),
    .io_ho_input(bc_pe_372_io_ho_input),
    .io_ve_input(bc_pe_372_io_ve_input),
    .io_input_valid(bc_pe_372_io_input_valid),
    .io_iormac(bc_pe_372_io_iormac),
    .io_ve_out(bc_pe_372_io_ve_out),
    .io_ho_out(bc_pe_372_io_ho_out),
    .io_res_out(bc_pe_372_io_res_out)
  );
  bc_pe bc_pe_373 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_373_clock),
    .reset(bc_pe_373_reset),
    .io_ho_input(bc_pe_373_io_ho_input),
    .io_ve_input(bc_pe_373_io_ve_input),
    .io_input_valid(bc_pe_373_io_input_valid),
    .io_iormac(bc_pe_373_io_iormac),
    .io_ve_out(bc_pe_373_io_ve_out),
    .io_ho_out(bc_pe_373_io_ho_out),
    .io_res_out(bc_pe_373_io_res_out)
  );
  bc_pe bc_pe_374 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_374_clock),
    .reset(bc_pe_374_reset),
    .io_ho_input(bc_pe_374_io_ho_input),
    .io_ve_input(bc_pe_374_io_ve_input),
    .io_input_valid(bc_pe_374_io_input_valid),
    .io_iormac(bc_pe_374_io_iormac),
    .io_ve_out(bc_pe_374_io_ve_out),
    .io_ho_out(bc_pe_374_io_ho_out),
    .io_res_out(bc_pe_374_io_res_out)
  );
  bc_pe bc_pe_375 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_375_clock),
    .reset(bc_pe_375_reset),
    .io_ho_input(bc_pe_375_io_ho_input),
    .io_ve_input(bc_pe_375_io_ve_input),
    .io_input_valid(bc_pe_375_io_input_valid),
    .io_iormac(bc_pe_375_io_iormac),
    .io_ve_out(bc_pe_375_io_ve_out),
    .io_ho_out(bc_pe_375_io_ho_out),
    .io_res_out(bc_pe_375_io_res_out)
  );
  bc_pe bc_pe_376 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_376_clock),
    .reset(bc_pe_376_reset),
    .io_ho_input(bc_pe_376_io_ho_input),
    .io_ve_input(bc_pe_376_io_ve_input),
    .io_input_valid(bc_pe_376_io_input_valid),
    .io_iormac(bc_pe_376_io_iormac),
    .io_ve_out(bc_pe_376_io_ve_out),
    .io_ho_out(bc_pe_376_io_ho_out),
    .io_res_out(bc_pe_376_io_res_out)
  );
  bc_pe bc_pe_377 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_377_clock),
    .reset(bc_pe_377_reset),
    .io_ho_input(bc_pe_377_io_ho_input),
    .io_ve_input(bc_pe_377_io_ve_input),
    .io_input_valid(bc_pe_377_io_input_valid),
    .io_iormac(bc_pe_377_io_iormac),
    .io_ve_out(bc_pe_377_io_ve_out),
    .io_ho_out(bc_pe_377_io_ho_out),
    .io_res_out(bc_pe_377_io_res_out)
  );
  bc_pe bc_pe_378 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_378_clock),
    .reset(bc_pe_378_reset),
    .io_ho_input(bc_pe_378_io_ho_input),
    .io_ve_input(bc_pe_378_io_ve_input),
    .io_input_valid(bc_pe_378_io_input_valid),
    .io_iormac(bc_pe_378_io_iormac),
    .io_ve_out(bc_pe_378_io_ve_out),
    .io_ho_out(bc_pe_378_io_ho_out),
    .io_res_out(bc_pe_378_io_res_out)
  );
  bc_pe bc_pe_379 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_379_clock),
    .reset(bc_pe_379_reset),
    .io_ho_input(bc_pe_379_io_ho_input),
    .io_ve_input(bc_pe_379_io_ve_input),
    .io_input_valid(bc_pe_379_io_input_valid),
    .io_iormac(bc_pe_379_io_iormac),
    .io_ve_out(bc_pe_379_io_ve_out),
    .io_ho_out(bc_pe_379_io_ho_out),
    .io_res_out(bc_pe_379_io_res_out)
  );
  bc_pe bc_pe_380 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_380_clock),
    .reset(bc_pe_380_reset),
    .io_ho_input(bc_pe_380_io_ho_input),
    .io_ve_input(bc_pe_380_io_ve_input),
    .io_input_valid(bc_pe_380_io_input_valid),
    .io_iormac(bc_pe_380_io_iormac),
    .io_ve_out(bc_pe_380_io_ve_out),
    .io_ho_out(bc_pe_380_io_ho_out),
    .io_res_out(bc_pe_380_io_res_out)
  );
  bc_pe bc_pe_381 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_381_clock),
    .reset(bc_pe_381_reset),
    .io_ho_input(bc_pe_381_io_ho_input),
    .io_ve_input(bc_pe_381_io_ve_input),
    .io_input_valid(bc_pe_381_io_input_valid),
    .io_iormac(bc_pe_381_io_iormac),
    .io_ve_out(bc_pe_381_io_ve_out),
    .io_ho_out(bc_pe_381_io_ho_out),
    .io_res_out(bc_pe_381_io_res_out)
  );
  bc_pe bc_pe_382 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_382_clock),
    .reset(bc_pe_382_reset),
    .io_ho_input(bc_pe_382_io_ho_input),
    .io_ve_input(bc_pe_382_io_ve_input),
    .io_input_valid(bc_pe_382_io_input_valid),
    .io_iormac(bc_pe_382_io_iormac),
    .io_ve_out(bc_pe_382_io_ve_out),
    .io_ho_out(bc_pe_382_io_ho_out),
    .io_res_out(bc_pe_382_io_res_out)
  );
  bc_pe bc_pe_383 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_383_clock),
    .reset(bc_pe_383_reset),
    .io_ho_input(bc_pe_383_io_ho_input),
    .io_ve_input(bc_pe_383_io_ve_input),
    .io_input_valid(bc_pe_383_io_input_valid),
    .io_iormac(bc_pe_383_io_iormac),
    .io_ve_out(bc_pe_383_io_ve_out),
    .io_ho_out(bc_pe_383_io_ho_out),
    .io_res_out(bc_pe_383_io_res_out)
  );
  bc_pe bc_pe_384 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_384_clock),
    .reset(bc_pe_384_reset),
    .io_ho_input(bc_pe_384_io_ho_input),
    .io_ve_input(bc_pe_384_io_ve_input),
    .io_input_valid(bc_pe_384_io_input_valid),
    .io_iormac(bc_pe_384_io_iormac),
    .io_ve_out(bc_pe_384_io_ve_out),
    .io_ho_out(bc_pe_384_io_ho_out),
    .io_res_out(bc_pe_384_io_res_out)
  );
  bc_pe bc_pe_385 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_385_clock),
    .reset(bc_pe_385_reset),
    .io_ho_input(bc_pe_385_io_ho_input),
    .io_ve_input(bc_pe_385_io_ve_input),
    .io_input_valid(bc_pe_385_io_input_valid),
    .io_iormac(bc_pe_385_io_iormac),
    .io_ve_out(bc_pe_385_io_ve_out),
    .io_ho_out(bc_pe_385_io_ho_out),
    .io_res_out(bc_pe_385_io_res_out)
  );
  bc_pe bc_pe_386 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_386_clock),
    .reset(bc_pe_386_reset),
    .io_ho_input(bc_pe_386_io_ho_input),
    .io_ve_input(bc_pe_386_io_ve_input),
    .io_input_valid(bc_pe_386_io_input_valid),
    .io_iormac(bc_pe_386_io_iormac),
    .io_ve_out(bc_pe_386_io_ve_out),
    .io_ho_out(bc_pe_386_io_ho_out),
    .io_res_out(bc_pe_386_io_res_out)
  );
  bc_pe bc_pe_387 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_387_clock),
    .reset(bc_pe_387_reset),
    .io_ho_input(bc_pe_387_io_ho_input),
    .io_ve_input(bc_pe_387_io_ve_input),
    .io_input_valid(bc_pe_387_io_input_valid),
    .io_iormac(bc_pe_387_io_iormac),
    .io_ve_out(bc_pe_387_io_ve_out),
    .io_ho_out(bc_pe_387_io_ho_out),
    .io_res_out(bc_pe_387_io_res_out)
  );
  bc_pe bc_pe_388 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_388_clock),
    .reset(bc_pe_388_reset),
    .io_ho_input(bc_pe_388_io_ho_input),
    .io_ve_input(bc_pe_388_io_ve_input),
    .io_input_valid(bc_pe_388_io_input_valid),
    .io_iormac(bc_pe_388_io_iormac),
    .io_ve_out(bc_pe_388_io_ve_out),
    .io_ho_out(bc_pe_388_io_ho_out),
    .io_res_out(bc_pe_388_io_res_out)
  );
  bc_pe bc_pe_389 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_389_clock),
    .reset(bc_pe_389_reset),
    .io_ho_input(bc_pe_389_io_ho_input),
    .io_ve_input(bc_pe_389_io_ve_input),
    .io_input_valid(bc_pe_389_io_input_valid),
    .io_iormac(bc_pe_389_io_iormac),
    .io_ve_out(bc_pe_389_io_ve_out),
    .io_ho_out(bc_pe_389_io_ho_out),
    .io_res_out(bc_pe_389_io_res_out)
  );
  bc_pe bc_pe_390 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_390_clock),
    .reset(bc_pe_390_reset),
    .io_ho_input(bc_pe_390_io_ho_input),
    .io_ve_input(bc_pe_390_io_ve_input),
    .io_input_valid(bc_pe_390_io_input_valid),
    .io_iormac(bc_pe_390_io_iormac),
    .io_ve_out(bc_pe_390_io_ve_out),
    .io_ho_out(bc_pe_390_io_ho_out),
    .io_res_out(bc_pe_390_io_res_out)
  );
  bc_pe bc_pe_391 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_391_clock),
    .reset(bc_pe_391_reset),
    .io_ho_input(bc_pe_391_io_ho_input),
    .io_ve_input(bc_pe_391_io_ve_input),
    .io_input_valid(bc_pe_391_io_input_valid),
    .io_iormac(bc_pe_391_io_iormac),
    .io_ve_out(bc_pe_391_io_ve_out),
    .io_ho_out(bc_pe_391_io_ho_out),
    .io_res_out(bc_pe_391_io_res_out)
  );
  bc_pe bc_pe_392 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_392_clock),
    .reset(bc_pe_392_reset),
    .io_ho_input(bc_pe_392_io_ho_input),
    .io_ve_input(bc_pe_392_io_ve_input),
    .io_input_valid(bc_pe_392_io_input_valid),
    .io_iormac(bc_pe_392_io_iormac),
    .io_ve_out(bc_pe_392_io_ve_out),
    .io_ho_out(bc_pe_392_io_ho_out),
    .io_res_out(bc_pe_392_io_res_out)
  );
  bc_pe bc_pe_393 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_393_clock),
    .reset(bc_pe_393_reset),
    .io_ho_input(bc_pe_393_io_ho_input),
    .io_ve_input(bc_pe_393_io_ve_input),
    .io_input_valid(bc_pe_393_io_input_valid),
    .io_iormac(bc_pe_393_io_iormac),
    .io_ve_out(bc_pe_393_io_ve_out),
    .io_ho_out(bc_pe_393_io_ho_out),
    .io_res_out(bc_pe_393_io_res_out)
  );
  bc_pe bc_pe_394 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_394_clock),
    .reset(bc_pe_394_reset),
    .io_ho_input(bc_pe_394_io_ho_input),
    .io_ve_input(bc_pe_394_io_ve_input),
    .io_input_valid(bc_pe_394_io_input_valid),
    .io_iormac(bc_pe_394_io_iormac),
    .io_ve_out(bc_pe_394_io_ve_out),
    .io_ho_out(bc_pe_394_io_ho_out),
    .io_res_out(bc_pe_394_io_res_out)
  );
  bc_pe bc_pe_395 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_395_clock),
    .reset(bc_pe_395_reset),
    .io_ho_input(bc_pe_395_io_ho_input),
    .io_ve_input(bc_pe_395_io_ve_input),
    .io_input_valid(bc_pe_395_io_input_valid),
    .io_iormac(bc_pe_395_io_iormac),
    .io_ve_out(bc_pe_395_io_ve_out),
    .io_ho_out(bc_pe_395_io_ho_out),
    .io_res_out(bc_pe_395_io_res_out)
  );
  bc_pe bc_pe_396 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_396_clock),
    .reset(bc_pe_396_reset),
    .io_ho_input(bc_pe_396_io_ho_input),
    .io_ve_input(bc_pe_396_io_ve_input),
    .io_input_valid(bc_pe_396_io_input_valid),
    .io_iormac(bc_pe_396_io_iormac),
    .io_ve_out(bc_pe_396_io_ve_out),
    .io_ho_out(bc_pe_396_io_ho_out),
    .io_res_out(bc_pe_396_io_res_out)
  );
  bc_pe bc_pe_397 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_397_clock),
    .reset(bc_pe_397_reset),
    .io_ho_input(bc_pe_397_io_ho_input),
    .io_ve_input(bc_pe_397_io_ve_input),
    .io_input_valid(bc_pe_397_io_input_valid),
    .io_iormac(bc_pe_397_io_iormac),
    .io_ve_out(bc_pe_397_io_ve_out),
    .io_ho_out(bc_pe_397_io_ho_out),
    .io_res_out(bc_pe_397_io_res_out)
  );
  bc_pe bc_pe_398 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_398_clock),
    .reset(bc_pe_398_reset),
    .io_ho_input(bc_pe_398_io_ho_input),
    .io_ve_input(bc_pe_398_io_ve_input),
    .io_input_valid(bc_pe_398_io_input_valid),
    .io_iormac(bc_pe_398_io_iormac),
    .io_ve_out(bc_pe_398_io_ve_out),
    .io_ho_out(bc_pe_398_io_ho_out),
    .io_res_out(bc_pe_398_io_res_out)
  );
  bc_pe bc_pe_399 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_399_clock),
    .reset(bc_pe_399_reset),
    .io_ho_input(bc_pe_399_io_ho_input),
    .io_ve_input(bc_pe_399_io_ve_input),
    .io_input_valid(bc_pe_399_io_input_valid),
    .io_iormac(bc_pe_399_io_iormac),
    .io_ve_out(bc_pe_399_io_ve_out),
    .io_ho_out(bc_pe_399_io_ho_out),
    .io_res_out(bc_pe_399_io_res_out)
  );
  bc_pe bc_pe_400 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_400_clock),
    .reset(bc_pe_400_reset),
    .io_ho_input(bc_pe_400_io_ho_input),
    .io_ve_input(bc_pe_400_io_ve_input),
    .io_input_valid(bc_pe_400_io_input_valid),
    .io_iormac(bc_pe_400_io_iormac),
    .io_ve_out(bc_pe_400_io_ve_out),
    .io_ho_out(bc_pe_400_io_ho_out),
    .io_res_out(bc_pe_400_io_res_out)
  );
  bc_pe bc_pe_401 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_401_clock),
    .reset(bc_pe_401_reset),
    .io_ho_input(bc_pe_401_io_ho_input),
    .io_ve_input(bc_pe_401_io_ve_input),
    .io_input_valid(bc_pe_401_io_input_valid),
    .io_iormac(bc_pe_401_io_iormac),
    .io_ve_out(bc_pe_401_io_ve_out),
    .io_ho_out(bc_pe_401_io_ho_out),
    .io_res_out(bc_pe_401_io_res_out)
  );
  bc_pe bc_pe_402 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_402_clock),
    .reset(bc_pe_402_reset),
    .io_ho_input(bc_pe_402_io_ho_input),
    .io_ve_input(bc_pe_402_io_ve_input),
    .io_input_valid(bc_pe_402_io_input_valid),
    .io_iormac(bc_pe_402_io_iormac),
    .io_ve_out(bc_pe_402_io_ve_out),
    .io_ho_out(bc_pe_402_io_ho_out),
    .io_res_out(bc_pe_402_io_res_out)
  );
  bc_pe bc_pe_403 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_403_clock),
    .reset(bc_pe_403_reset),
    .io_ho_input(bc_pe_403_io_ho_input),
    .io_ve_input(bc_pe_403_io_ve_input),
    .io_input_valid(bc_pe_403_io_input_valid),
    .io_iormac(bc_pe_403_io_iormac),
    .io_ve_out(bc_pe_403_io_ve_out),
    .io_ho_out(bc_pe_403_io_ho_out),
    .io_res_out(bc_pe_403_io_res_out)
  );
  bc_pe bc_pe_404 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_404_clock),
    .reset(bc_pe_404_reset),
    .io_ho_input(bc_pe_404_io_ho_input),
    .io_ve_input(bc_pe_404_io_ve_input),
    .io_input_valid(bc_pe_404_io_input_valid),
    .io_iormac(bc_pe_404_io_iormac),
    .io_ve_out(bc_pe_404_io_ve_out),
    .io_ho_out(bc_pe_404_io_ho_out),
    .io_res_out(bc_pe_404_io_res_out)
  );
  bc_pe bc_pe_405 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_405_clock),
    .reset(bc_pe_405_reset),
    .io_ho_input(bc_pe_405_io_ho_input),
    .io_ve_input(bc_pe_405_io_ve_input),
    .io_input_valid(bc_pe_405_io_input_valid),
    .io_iormac(bc_pe_405_io_iormac),
    .io_ve_out(bc_pe_405_io_ve_out),
    .io_ho_out(bc_pe_405_io_ho_out),
    .io_res_out(bc_pe_405_io_res_out)
  );
  bc_pe bc_pe_406 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_406_clock),
    .reset(bc_pe_406_reset),
    .io_ho_input(bc_pe_406_io_ho_input),
    .io_ve_input(bc_pe_406_io_ve_input),
    .io_input_valid(bc_pe_406_io_input_valid),
    .io_iormac(bc_pe_406_io_iormac),
    .io_ve_out(bc_pe_406_io_ve_out),
    .io_ho_out(bc_pe_406_io_ho_out),
    .io_res_out(bc_pe_406_io_res_out)
  );
  bc_pe bc_pe_407 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_407_clock),
    .reset(bc_pe_407_reset),
    .io_ho_input(bc_pe_407_io_ho_input),
    .io_ve_input(bc_pe_407_io_ve_input),
    .io_input_valid(bc_pe_407_io_input_valid),
    .io_iormac(bc_pe_407_io_iormac),
    .io_ve_out(bc_pe_407_io_ve_out),
    .io_ho_out(bc_pe_407_io_ho_out),
    .io_res_out(bc_pe_407_io_res_out)
  );
  bc_pe bc_pe_408 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_408_clock),
    .reset(bc_pe_408_reset),
    .io_ho_input(bc_pe_408_io_ho_input),
    .io_ve_input(bc_pe_408_io_ve_input),
    .io_input_valid(bc_pe_408_io_input_valid),
    .io_iormac(bc_pe_408_io_iormac),
    .io_ve_out(bc_pe_408_io_ve_out),
    .io_ho_out(bc_pe_408_io_ho_out),
    .io_res_out(bc_pe_408_io_res_out)
  );
  bc_pe bc_pe_409 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_409_clock),
    .reset(bc_pe_409_reset),
    .io_ho_input(bc_pe_409_io_ho_input),
    .io_ve_input(bc_pe_409_io_ve_input),
    .io_input_valid(bc_pe_409_io_input_valid),
    .io_iormac(bc_pe_409_io_iormac),
    .io_ve_out(bc_pe_409_io_ve_out),
    .io_ho_out(bc_pe_409_io_ho_out),
    .io_res_out(bc_pe_409_io_res_out)
  );
  bc_pe bc_pe_410 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_410_clock),
    .reset(bc_pe_410_reset),
    .io_ho_input(bc_pe_410_io_ho_input),
    .io_ve_input(bc_pe_410_io_ve_input),
    .io_input_valid(bc_pe_410_io_input_valid),
    .io_iormac(bc_pe_410_io_iormac),
    .io_ve_out(bc_pe_410_io_ve_out),
    .io_ho_out(bc_pe_410_io_ho_out),
    .io_res_out(bc_pe_410_io_res_out)
  );
  bc_pe bc_pe_411 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_411_clock),
    .reset(bc_pe_411_reset),
    .io_ho_input(bc_pe_411_io_ho_input),
    .io_ve_input(bc_pe_411_io_ve_input),
    .io_input_valid(bc_pe_411_io_input_valid),
    .io_iormac(bc_pe_411_io_iormac),
    .io_ve_out(bc_pe_411_io_ve_out),
    .io_ho_out(bc_pe_411_io_ho_out),
    .io_res_out(bc_pe_411_io_res_out)
  );
  bc_pe bc_pe_412 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_412_clock),
    .reset(bc_pe_412_reset),
    .io_ho_input(bc_pe_412_io_ho_input),
    .io_ve_input(bc_pe_412_io_ve_input),
    .io_input_valid(bc_pe_412_io_input_valid),
    .io_iormac(bc_pe_412_io_iormac),
    .io_ve_out(bc_pe_412_io_ve_out),
    .io_ho_out(bc_pe_412_io_ho_out),
    .io_res_out(bc_pe_412_io_res_out)
  );
  bc_pe bc_pe_413 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_413_clock),
    .reset(bc_pe_413_reset),
    .io_ho_input(bc_pe_413_io_ho_input),
    .io_ve_input(bc_pe_413_io_ve_input),
    .io_input_valid(bc_pe_413_io_input_valid),
    .io_iormac(bc_pe_413_io_iormac),
    .io_ve_out(bc_pe_413_io_ve_out),
    .io_ho_out(bc_pe_413_io_ho_out),
    .io_res_out(bc_pe_413_io_res_out)
  );
  bc_pe bc_pe_414 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_414_clock),
    .reset(bc_pe_414_reset),
    .io_ho_input(bc_pe_414_io_ho_input),
    .io_ve_input(bc_pe_414_io_ve_input),
    .io_input_valid(bc_pe_414_io_input_valid),
    .io_iormac(bc_pe_414_io_iormac),
    .io_ve_out(bc_pe_414_io_ve_out),
    .io_ho_out(bc_pe_414_io_ho_out),
    .io_res_out(bc_pe_414_io_res_out)
  );
  bc_pe bc_pe_415 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_415_clock),
    .reset(bc_pe_415_reset),
    .io_ho_input(bc_pe_415_io_ho_input),
    .io_ve_input(bc_pe_415_io_ve_input),
    .io_input_valid(bc_pe_415_io_input_valid),
    .io_iormac(bc_pe_415_io_iormac),
    .io_ve_out(bc_pe_415_io_ve_out),
    .io_ho_out(bc_pe_415_io_ho_out),
    .io_res_out(bc_pe_415_io_res_out)
  );
  bc_pe bc_pe_416 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_416_clock),
    .reset(bc_pe_416_reset),
    .io_ho_input(bc_pe_416_io_ho_input),
    .io_ve_input(bc_pe_416_io_ve_input),
    .io_input_valid(bc_pe_416_io_input_valid),
    .io_iormac(bc_pe_416_io_iormac),
    .io_ve_out(bc_pe_416_io_ve_out),
    .io_ho_out(bc_pe_416_io_ho_out),
    .io_res_out(bc_pe_416_io_res_out)
  );
  bc_pe bc_pe_417 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_417_clock),
    .reset(bc_pe_417_reset),
    .io_ho_input(bc_pe_417_io_ho_input),
    .io_ve_input(bc_pe_417_io_ve_input),
    .io_input_valid(bc_pe_417_io_input_valid),
    .io_iormac(bc_pe_417_io_iormac),
    .io_ve_out(bc_pe_417_io_ve_out),
    .io_ho_out(bc_pe_417_io_ho_out),
    .io_res_out(bc_pe_417_io_res_out)
  );
  bc_pe bc_pe_418 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_418_clock),
    .reset(bc_pe_418_reset),
    .io_ho_input(bc_pe_418_io_ho_input),
    .io_ve_input(bc_pe_418_io_ve_input),
    .io_input_valid(bc_pe_418_io_input_valid),
    .io_iormac(bc_pe_418_io_iormac),
    .io_ve_out(bc_pe_418_io_ve_out),
    .io_ho_out(bc_pe_418_io_ho_out),
    .io_res_out(bc_pe_418_io_res_out)
  );
  bc_pe bc_pe_419 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_419_clock),
    .reset(bc_pe_419_reset),
    .io_ho_input(bc_pe_419_io_ho_input),
    .io_ve_input(bc_pe_419_io_ve_input),
    .io_input_valid(bc_pe_419_io_input_valid),
    .io_iormac(bc_pe_419_io_iormac),
    .io_ve_out(bc_pe_419_io_ve_out),
    .io_ho_out(bc_pe_419_io_ho_out),
    .io_res_out(bc_pe_419_io_res_out)
  );
  bc_pe bc_pe_420 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_420_clock),
    .reset(bc_pe_420_reset),
    .io_ho_input(bc_pe_420_io_ho_input),
    .io_ve_input(bc_pe_420_io_ve_input),
    .io_input_valid(bc_pe_420_io_input_valid),
    .io_iormac(bc_pe_420_io_iormac),
    .io_ve_out(bc_pe_420_io_ve_out),
    .io_ho_out(bc_pe_420_io_ho_out),
    .io_res_out(bc_pe_420_io_res_out)
  );
  bc_pe bc_pe_421 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_421_clock),
    .reset(bc_pe_421_reset),
    .io_ho_input(bc_pe_421_io_ho_input),
    .io_ve_input(bc_pe_421_io_ve_input),
    .io_input_valid(bc_pe_421_io_input_valid),
    .io_iormac(bc_pe_421_io_iormac),
    .io_ve_out(bc_pe_421_io_ve_out),
    .io_ho_out(bc_pe_421_io_ho_out),
    .io_res_out(bc_pe_421_io_res_out)
  );
  bc_pe bc_pe_422 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_422_clock),
    .reset(bc_pe_422_reset),
    .io_ho_input(bc_pe_422_io_ho_input),
    .io_ve_input(bc_pe_422_io_ve_input),
    .io_input_valid(bc_pe_422_io_input_valid),
    .io_iormac(bc_pe_422_io_iormac),
    .io_ve_out(bc_pe_422_io_ve_out),
    .io_ho_out(bc_pe_422_io_ho_out),
    .io_res_out(bc_pe_422_io_res_out)
  );
  bc_pe bc_pe_423 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_423_clock),
    .reset(bc_pe_423_reset),
    .io_ho_input(bc_pe_423_io_ho_input),
    .io_ve_input(bc_pe_423_io_ve_input),
    .io_input_valid(bc_pe_423_io_input_valid),
    .io_iormac(bc_pe_423_io_iormac),
    .io_ve_out(bc_pe_423_io_ve_out),
    .io_ho_out(bc_pe_423_io_ho_out),
    .io_res_out(bc_pe_423_io_res_out)
  );
  bc_pe bc_pe_424 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_424_clock),
    .reset(bc_pe_424_reset),
    .io_ho_input(bc_pe_424_io_ho_input),
    .io_ve_input(bc_pe_424_io_ve_input),
    .io_input_valid(bc_pe_424_io_input_valid),
    .io_iormac(bc_pe_424_io_iormac),
    .io_ve_out(bc_pe_424_io_ve_out),
    .io_ho_out(bc_pe_424_io_ho_out),
    .io_res_out(bc_pe_424_io_res_out)
  );
  bc_pe bc_pe_425 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_425_clock),
    .reset(bc_pe_425_reset),
    .io_ho_input(bc_pe_425_io_ho_input),
    .io_ve_input(bc_pe_425_io_ve_input),
    .io_input_valid(bc_pe_425_io_input_valid),
    .io_iormac(bc_pe_425_io_iormac),
    .io_ve_out(bc_pe_425_io_ve_out),
    .io_ho_out(bc_pe_425_io_ho_out),
    .io_res_out(bc_pe_425_io_res_out)
  );
  bc_pe bc_pe_426 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_426_clock),
    .reset(bc_pe_426_reset),
    .io_ho_input(bc_pe_426_io_ho_input),
    .io_ve_input(bc_pe_426_io_ve_input),
    .io_input_valid(bc_pe_426_io_input_valid),
    .io_iormac(bc_pe_426_io_iormac),
    .io_ve_out(bc_pe_426_io_ve_out),
    .io_ho_out(bc_pe_426_io_ho_out),
    .io_res_out(bc_pe_426_io_res_out)
  );
  bc_pe bc_pe_427 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_427_clock),
    .reset(bc_pe_427_reset),
    .io_ho_input(bc_pe_427_io_ho_input),
    .io_ve_input(bc_pe_427_io_ve_input),
    .io_input_valid(bc_pe_427_io_input_valid),
    .io_iormac(bc_pe_427_io_iormac),
    .io_ve_out(bc_pe_427_io_ve_out),
    .io_ho_out(bc_pe_427_io_ho_out),
    .io_res_out(bc_pe_427_io_res_out)
  );
  bc_pe bc_pe_428 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_428_clock),
    .reset(bc_pe_428_reset),
    .io_ho_input(bc_pe_428_io_ho_input),
    .io_ve_input(bc_pe_428_io_ve_input),
    .io_input_valid(bc_pe_428_io_input_valid),
    .io_iormac(bc_pe_428_io_iormac),
    .io_ve_out(bc_pe_428_io_ve_out),
    .io_ho_out(bc_pe_428_io_ho_out),
    .io_res_out(bc_pe_428_io_res_out)
  );
  bc_pe bc_pe_429 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_429_clock),
    .reset(bc_pe_429_reset),
    .io_ho_input(bc_pe_429_io_ho_input),
    .io_ve_input(bc_pe_429_io_ve_input),
    .io_input_valid(bc_pe_429_io_input_valid),
    .io_iormac(bc_pe_429_io_iormac),
    .io_ve_out(bc_pe_429_io_ve_out),
    .io_ho_out(bc_pe_429_io_ho_out),
    .io_res_out(bc_pe_429_io_res_out)
  );
  bc_pe bc_pe_430 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_430_clock),
    .reset(bc_pe_430_reset),
    .io_ho_input(bc_pe_430_io_ho_input),
    .io_ve_input(bc_pe_430_io_ve_input),
    .io_input_valid(bc_pe_430_io_input_valid),
    .io_iormac(bc_pe_430_io_iormac),
    .io_ve_out(bc_pe_430_io_ve_out),
    .io_ho_out(bc_pe_430_io_ho_out),
    .io_res_out(bc_pe_430_io_res_out)
  );
  bc_pe bc_pe_431 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_431_clock),
    .reset(bc_pe_431_reset),
    .io_ho_input(bc_pe_431_io_ho_input),
    .io_ve_input(bc_pe_431_io_ve_input),
    .io_input_valid(bc_pe_431_io_input_valid),
    .io_iormac(bc_pe_431_io_iormac),
    .io_ve_out(bc_pe_431_io_ve_out),
    .io_ho_out(bc_pe_431_io_ho_out),
    .io_res_out(bc_pe_431_io_res_out)
  );
  bc_pe bc_pe_432 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_432_clock),
    .reset(bc_pe_432_reset),
    .io_ho_input(bc_pe_432_io_ho_input),
    .io_ve_input(bc_pe_432_io_ve_input),
    .io_input_valid(bc_pe_432_io_input_valid),
    .io_iormac(bc_pe_432_io_iormac),
    .io_ve_out(bc_pe_432_io_ve_out),
    .io_ho_out(bc_pe_432_io_ho_out),
    .io_res_out(bc_pe_432_io_res_out)
  );
  bc_pe bc_pe_433 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_433_clock),
    .reset(bc_pe_433_reset),
    .io_ho_input(bc_pe_433_io_ho_input),
    .io_ve_input(bc_pe_433_io_ve_input),
    .io_input_valid(bc_pe_433_io_input_valid),
    .io_iormac(bc_pe_433_io_iormac),
    .io_ve_out(bc_pe_433_io_ve_out),
    .io_ho_out(bc_pe_433_io_ho_out),
    .io_res_out(bc_pe_433_io_res_out)
  );
  bc_pe bc_pe_434 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_434_clock),
    .reset(bc_pe_434_reset),
    .io_ho_input(bc_pe_434_io_ho_input),
    .io_ve_input(bc_pe_434_io_ve_input),
    .io_input_valid(bc_pe_434_io_input_valid),
    .io_iormac(bc_pe_434_io_iormac),
    .io_ve_out(bc_pe_434_io_ve_out),
    .io_ho_out(bc_pe_434_io_ho_out),
    .io_res_out(bc_pe_434_io_res_out)
  );
  bc_pe bc_pe_435 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_435_clock),
    .reset(bc_pe_435_reset),
    .io_ho_input(bc_pe_435_io_ho_input),
    .io_ve_input(bc_pe_435_io_ve_input),
    .io_input_valid(bc_pe_435_io_input_valid),
    .io_iormac(bc_pe_435_io_iormac),
    .io_ve_out(bc_pe_435_io_ve_out),
    .io_ho_out(bc_pe_435_io_ho_out),
    .io_res_out(bc_pe_435_io_res_out)
  );
  bc_pe bc_pe_436 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_436_clock),
    .reset(bc_pe_436_reset),
    .io_ho_input(bc_pe_436_io_ho_input),
    .io_ve_input(bc_pe_436_io_ve_input),
    .io_input_valid(bc_pe_436_io_input_valid),
    .io_iormac(bc_pe_436_io_iormac),
    .io_ve_out(bc_pe_436_io_ve_out),
    .io_ho_out(bc_pe_436_io_ho_out),
    .io_res_out(bc_pe_436_io_res_out)
  );
  bc_pe bc_pe_437 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_437_clock),
    .reset(bc_pe_437_reset),
    .io_ho_input(bc_pe_437_io_ho_input),
    .io_ve_input(bc_pe_437_io_ve_input),
    .io_input_valid(bc_pe_437_io_input_valid),
    .io_iormac(bc_pe_437_io_iormac),
    .io_ve_out(bc_pe_437_io_ve_out),
    .io_ho_out(bc_pe_437_io_ho_out),
    .io_res_out(bc_pe_437_io_res_out)
  );
  bc_pe bc_pe_438 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_438_clock),
    .reset(bc_pe_438_reset),
    .io_ho_input(bc_pe_438_io_ho_input),
    .io_ve_input(bc_pe_438_io_ve_input),
    .io_input_valid(bc_pe_438_io_input_valid),
    .io_iormac(bc_pe_438_io_iormac),
    .io_ve_out(bc_pe_438_io_ve_out),
    .io_ho_out(bc_pe_438_io_ho_out),
    .io_res_out(bc_pe_438_io_res_out)
  );
  bc_pe bc_pe_439 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_439_clock),
    .reset(bc_pe_439_reset),
    .io_ho_input(bc_pe_439_io_ho_input),
    .io_ve_input(bc_pe_439_io_ve_input),
    .io_input_valid(bc_pe_439_io_input_valid),
    .io_iormac(bc_pe_439_io_iormac),
    .io_ve_out(bc_pe_439_io_ve_out),
    .io_ho_out(bc_pe_439_io_ho_out),
    .io_res_out(bc_pe_439_io_res_out)
  );
  bc_pe bc_pe_440 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_440_clock),
    .reset(bc_pe_440_reset),
    .io_ho_input(bc_pe_440_io_ho_input),
    .io_ve_input(bc_pe_440_io_ve_input),
    .io_input_valid(bc_pe_440_io_input_valid),
    .io_iormac(bc_pe_440_io_iormac),
    .io_ve_out(bc_pe_440_io_ve_out),
    .io_ho_out(bc_pe_440_io_ho_out),
    .io_res_out(bc_pe_440_io_res_out)
  );
  bc_pe bc_pe_441 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_441_clock),
    .reset(bc_pe_441_reset),
    .io_ho_input(bc_pe_441_io_ho_input),
    .io_ve_input(bc_pe_441_io_ve_input),
    .io_input_valid(bc_pe_441_io_input_valid),
    .io_iormac(bc_pe_441_io_iormac),
    .io_ve_out(bc_pe_441_io_ve_out),
    .io_ho_out(bc_pe_441_io_ho_out),
    .io_res_out(bc_pe_441_io_res_out)
  );
  bc_pe bc_pe_442 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_442_clock),
    .reset(bc_pe_442_reset),
    .io_ho_input(bc_pe_442_io_ho_input),
    .io_ve_input(bc_pe_442_io_ve_input),
    .io_input_valid(bc_pe_442_io_input_valid),
    .io_iormac(bc_pe_442_io_iormac),
    .io_ve_out(bc_pe_442_io_ve_out),
    .io_ho_out(bc_pe_442_io_ho_out),
    .io_res_out(bc_pe_442_io_res_out)
  );
  bc_pe bc_pe_443 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_443_clock),
    .reset(bc_pe_443_reset),
    .io_ho_input(bc_pe_443_io_ho_input),
    .io_ve_input(bc_pe_443_io_ve_input),
    .io_input_valid(bc_pe_443_io_input_valid),
    .io_iormac(bc_pe_443_io_iormac),
    .io_ve_out(bc_pe_443_io_ve_out),
    .io_ho_out(bc_pe_443_io_ho_out),
    .io_res_out(bc_pe_443_io_res_out)
  );
  bc_pe bc_pe_444 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_444_clock),
    .reset(bc_pe_444_reset),
    .io_ho_input(bc_pe_444_io_ho_input),
    .io_ve_input(bc_pe_444_io_ve_input),
    .io_input_valid(bc_pe_444_io_input_valid),
    .io_iormac(bc_pe_444_io_iormac),
    .io_ve_out(bc_pe_444_io_ve_out),
    .io_ho_out(bc_pe_444_io_ho_out),
    .io_res_out(bc_pe_444_io_res_out)
  );
  bc_pe bc_pe_445 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_445_clock),
    .reset(bc_pe_445_reset),
    .io_ho_input(bc_pe_445_io_ho_input),
    .io_ve_input(bc_pe_445_io_ve_input),
    .io_input_valid(bc_pe_445_io_input_valid),
    .io_iormac(bc_pe_445_io_iormac),
    .io_ve_out(bc_pe_445_io_ve_out),
    .io_ho_out(bc_pe_445_io_ho_out),
    .io_res_out(bc_pe_445_io_res_out)
  );
  bc_pe bc_pe_446 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_446_clock),
    .reset(bc_pe_446_reset),
    .io_ho_input(bc_pe_446_io_ho_input),
    .io_ve_input(bc_pe_446_io_ve_input),
    .io_input_valid(bc_pe_446_io_input_valid),
    .io_iormac(bc_pe_446_io_iormac),
    .io_ve_out(bc_pe_446_io_ve_out),
    .io_ho_out(bc_pe_446_io_ho_out),
    .io_res_out(bc_pe_446_io_res_out)
  );
  bc_pe bc_pe_447 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_447_clock),
    .reset(bc_pe_447_reset),
    .io_ho_input(bc_pe_447_io_ho_input),
    .io_ve_input(bc_pe_447_io_ve_input),
    .io_input_valid(bc_pe_447_io_input_valid),
    .io_iormac(bc_pe_447_io_iormac),
    .io_ve_out(bc_pe_447_io_ve_out),
    .io_ho_out(bc_pe_447_io_ho_out),
    .io_res_out(bc_pe_447_io_res_out)
  );
  bc_pe bc_pe_448 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_448_clock),
    .reset(bc_pe_448_reset),
    .io_ho_input(bc_pe_448_io_ho_input),
    .io_ve_input(bc_pe_448_io_ve_input),
    .io_input_valid(bc_pe_448_io_input_valid),
    .io_iormac(bc_pe_448_io_iormac),
    .io_ve_out(bc_pe_448_io_ve_out),
    .io_ho_out(bc_pe_448_io_ho_out),
    .io_res_out(bc_pe_448_io_res_out)
  );
  bc_pe bc_pe_449 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_449_clock),
    .reset(bc_pe_449_reset),
    .io_ho_input(bc_pe_449_io_ho_input),
    .io_ve_input(bc_pe_449_io_ve_input),
    .io_input_valid(bc_pe_449_io_input_valid),
    .io_iormac(bc_pe_449_io_iormac),
    .io_ve_out(bc_pe_449_io_ve_out),
    .io_ho_out(bc_pe_449_io_ho_out),
    .io_res_out(bc_pe_449_io_res_out)
  );
  bc_pe bc_pe_450 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_450_clock),
    .reset(bc_pe_450_reset),
    .io_ho_input(bc_pe_450_io_ho_input),
    .io_ve_input(bc_pe_450_io_ve_input),
    .io_input_valid(bc_pe_450_io_input_valid),
    .io_iormac(bc_pe_450_io_iormac),
    .io_ve_out(bc_pe_450_io_ve_out),
    .io_ho_out(bc_pe_450_io_ho_out),
    .io_res_out(bc_pe_450_io_res_out)
  );
  bc_pe bc_pe_451 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_451_clock),
    .reset(bc_pe_451_reset),
    .io_ho_input(bc_pe_451_io_ho_input),
    .io_ve_input(bc_pe_451_io_ve_input),
    .io_input_valid(bc_pe_451_io_input_valid),
    .io_iormac(bc_pe_451_io_iormac),
    .io_ve_out(bc_pe_451_io_ve_out),
    .io_ho_out(bc_pe_451_io_ho_out),
    .io_res_out(bc_pe_451_io_res_out)
  );
  bc_pe bc_pe_452 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_452_clock),
    .reset(bc_pe_452_reset),
    .io_ho_input(bc_pe_452_io_ho_input),
    .io_ve_input(bc_pe_452_io_ve_input),
    .io_input_valid(bc_pe_452_io_input_valid),
    .io_iormac(bc_pe_452_io_iormac),
    .io_ve_out(bc_pe_452_io_ve_out),
    .io_ho_out(bc_pe_452_io_ho_out),
    .io_res_out(bc_pe_452_io_res_out)
  );
  bc_pe bc_pe_453 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_453_clock),
    .reset(bc_pe_453_reset),
    .io_ho_input(bc_pe_453_io_ho_input),
    .io_ve_input(bc_pe_453_io_ve_input),
    .io_input_valid(bc_pe_453_io_input_valid),
    .io_iormac(bc_pe_453_io_iormac),
    .io_ve_out(bc_pe_453_io_ve_out),
    .io_ho_out(bc_pe_453_io_ho_out),
    .io_res_out(bc_pe_453_io_res_out)
  );
  bc_pe bc_pe_454 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_454_clock),
    .reset(bc_pe_454_reset),
    .io_ho_input(bc_pe_454_io_ho_input),
    .io_ve_input(bc_pe_454_io_ve_input),
    .io_input_valid(bc_pe_454_io_input_valid),
    .io_iormac(bc_pe_454_io_iormac),
    .io_ve_out(bc_pe_454_io_ve_out),
    .io_ho_out(bc_pe_454_io_ho_out),
    .io_res_out(bc_pe_454_io_res_out)
  );
  bc_pe bc_pe_455 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_455_clock),
    .reset(bc_pe_455_reset),
    .io_ho_input(bc_pe_455_io_ho_input),
    .io_ve_input(bc_pe_455_io_ve_input),
    .io_input_valid(bc_pe_455_io_input_valid),
    .io_iormac(bc_pe_455_io_iormac),
    .io_ve_out(bc_pe_455_io_ve_out),
    .io_ho_out(bc_pe_455_io_ho_out),
    .io_res_out(bc_pe_455_io_res_out)
  );
  bc_pe bc_pe_456 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_456_clock),
    .reset(bc_pe_456_reset),
    .io_ho_input(bc_pe_456_io_ho_input),
    .io_ve_input(bc_pe_456_io_ve_input),
    .io_input_valid(bc_pe_456_io_input_valid),
    .io_iormac(bc_pe_456_io_iormac),
    .io_ve_out(bc_pe_456_io_ve_out),
    .io_ho_out(bc_pe_456_io_ho_out),
    .io_res_out(bc_pe_456_io_res_out)
  );
  bc_pe bc_pe_457 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_457_clock),
    .reset(bc_pe_457_reset),
    .io_ho_input(bc_pe_457_io_ho_input),
    .io_ve_input(bc_pe_457_io_ve_input),
    .io_input_valid(bc_pe_457_io_input_valid),
    .io_iormac(bc_pe_457_io_iormac),
    .io_ve_out(bc_pe_457_io_ve_out),
    .io_ho_out(bc_pe_457_io_ho_out),
    .io_res_out(bc_pe_457_io_res_out)
  );
  bc_pe bc_pe_458 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_458_clock),
    .reset(bc_pe_458_reset),
    .io_ho_input(bc_pe_458_io_ho_input),
    .io_ve_input(bc_pe_458_io_ve_input),
    .io_input_valid(bc_pe_458_io_input_valid),
    .io_iormac(bc_pe_458_io_iormac),
    .io_ve_out(bc_pe_458_io_ve_out),
    .io_ho_out(bc_pe_458_io_ho_out),
    .io_res_out(bc_pe_458_io_res_out)
  );
  bc_pe bc_pe_459 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_459_clock),
    .reset(bc_pe_459_reset),
    .io_ho_input(bc_pe_459_io_ho_input),
    .io_ve_input(bc_pe_459_io_ve_input),
    .io_input_valid(bc_pe_459_io_input_valid),
    .io_iormac(bc_pe_459_io_iormac),
    .io_ve_out(bc_pe_459_io_ve_out),
    .io_ho_out(bc_pe_459_io_ho_out),
    .io_res_out(bc_pe_459_io_res_out)
  );
  bc_pe bc_pe_460 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_460_clock),
    .reset(bc_pe_460_reset),
    .io_ho_input(bc_pe_460_io_ho_input),
    .io_ve_input(bc_pe_460_io_ve_input),
    .io_input_valid(bc_pe_460_io_input_valid),
    .io_iormac(bc_pe_460_io_iormac),
    .io_ve_out(bc_pe_460_io_ve_out),
    .io_ho_out(bc_pe_460_io_ho_out),
    .io_res_out(bc_pe_460_io_res_out)
  );
  bc_pe bc_pe_461 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_461_clock),
    .reset(bc_pe_461_reset),
    .io_ho_input(bc_pe_461_io_ho_input),
    .io_ve_input(bc_pe_461_io_ve_input),
    .io_input_valid(bc_pe_461_io_input_valid),
    .io_iormac(bc_pe_461_io_iormac),
    .io_ve_out(bc_pe_461_io_ve_out),
    .io_ho_out(bc_pe_461_io_ho_out),
    .io_res_out(bc_pe_461_io_res_out)
  );
  bc_pe bc_pe_462 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_462_clock),
    .reset(bc_pe_462_reset),
    .io_ho_input(bc_pe_462_io_ho_input),
    .io_ve_input(bc_pe_462_io_ve_input),
    .io_input_valid(bc_pe_462_io_input_valid),
    .io_iormac(bc_pe_462_io_iormac),
    .io_ve_out(bc_pe_462_io_ve_out),
    .io_ho_out(bc_pe_462_io_ho_out),
    .io_res_out(bc_pe_462_io_res_out)
  );
  bc_pe bc_pe_463 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_463_clock),
    .reset(bc_pe_463_reset),
    .io_ho_input(bc_pe_463_io_ho_input),
    .io_ve_input(bc_pe_463_io_ve_input),
    .io_input_valid(bc_pe_463_io_input_valid),
    .io_iormac(bc_pe_463_io_iormac),
    .io_ve_out(bc_pe_463_io_ve_out),
    .io_ho_out(bc_pe_463_io_ho_out),
    .io_res_out(bc_pe_463_io_res_out)
  );
  bc_pe bc_pe_464 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_464_clock),
    .reset(bc_pe_464_reset),
    .io_ho_input(bc_pe_464_io_ho_input),
    .io_ve_input(bc_pe_464_io_ve_input),
    .io_input_valid(bc_pe_464_io_input_valid),
    .io_iormac(bc_pe_464_io_iormac),
    .io_ve_out(bc_pe_464_io_ve_out),
    .io_ho_out(bc_pe_464_io_ho_out),
    .io_res_out(bc_pe_464_io_res_out)
  );
  bc_pe bc_pe_465 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_465_clock),
    .reset(bc_pe_465_reset),
    .io_ho_input(bc_pe_465_io_ho_input),
    .io_ve_input(bc_pe_465_io_ve_input),
    .io_input_valid(bc_pe_465_io_input_valid),
    .io_iormac(bc_pe_465_io_iormac),
    .io_ve_out(bc_pe_465_io_ve_out),
    .io_ho_out(bc_pe_465_io_ho_out),
    .io_res_out(bc_pe_465_io_res_out)
  );
  bc_pe bc_pe_466 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_466_clock),
    .reset(bc_pe_466_reset),
    .io_ho_input(bc_pe_466_io_ho_input),
    .io_ve_input(bc_pe_466_io_ve_input),
    .io_input_valid(bc_pe_466_io_input_valid),
    .io_iormac(bc_pe_466_io_iormac),
    .io_ve_out(bc_pe_466_io_ve_out),
    .io_ho_out(bc_pe_466_io_ho_out),
    .io_res_out(bc_pe_466_io_res_out)
  );
  bc_pe bc_pe_467 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_467_clock),
    .reset(bc_pe_467_reset),
    .io_ho_input(bc_pe_467_io_ho_input),
    .io_ve_input(bc_pe_467_io_ve_input),
    .io_input_valid(bc_pe_467_io_input_valid),
    .io_iormac(bc_pe_467_io_iormac),
    .io_ve_out(bc_pe_467_io_ve_out),
    .io_ho_out(bc_pe_467_io_ho_out),
    .io_res_out(bc_pe_467_io_res_out)
  );
  bc_pe bc_pe_468 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_468_clock),
    .reset(bc_pe_468_reset),
    .io_ho_input(bc_pe_468_io_ho_input),
    .io_ve_input(bc_pe_468_io_ve_input),
    .io_input_valid(bc_pe_468_io_input_valid),
    .io_iormac(bc_pe_468_io_iormac),
    .io_ve_out(bc_pe_468_io_ve_out),
    .io_ho_out(bc_pe_468_io_ho_out),
    .io_res_out(bc_pe_468_io_res_out)
  );
  bc_pe bc_pe_469 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_469_clock),
    .reset(bc_pe_469_reset),
    .io_ho_input(bc_pe_469_io_ho_input),
    .io_ve_input(bc_pe_469_io_ve_input),
    .io_input_valid(bc_pe_469_io_input_valid),
    .io_iormac(bc_pe_469_io_iormac),
    .io_ve_out(bc_pe_469_io_ve_out),
    .io_ho_out(bc_pe_469_io_ho_out),
    .io_res_out(bc_pe_469_io_res_out)
  );
  bc_pe bc_pe_470 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_470_clock),
    .reset(bc_pe_470_reset),
    .io_ho_input(bc_pe_470_io_ho_input),
    .io_ve_input(bc_pe_470_io_ve_input),
    .io_input_valid(bc_pe_470_io_input_valid),
    .io_iormac(bc_pe_470_io_iormac),
    .io_ve_out(bc_pe_470_io_ve_out),
    .io_ho_out(bc_pe_470_io_ho_out),
    .io_res_out(bc_pe_470_io_res_out)
  );
  bc_pe bc_pe_471 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_471_clock),
    .reset(bc_pe_471_reset),
    .io_ho_input(bc_pe_471_io_ho_input),
    .io_ve_input(bc_pe_471_io_ve_input),
    .io_input_valid(bc_pe_471_io_input_valid),
    .io_iormac(bc_pe_471_io_iormac),
    .io_ve_out(bc_pe_471_io_ve_out),
    .io_ho_out(bc_pe_471_io_ho_out),
    .io_res_out(bc_pe_471_io_res_out)
  );
  bc_pe bc_pe_472 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_472_clock),
    .reset(bc_pe_472_reset),
    .io_ho_input(bc_pe_472_io_ho_input),
    .io_ve_input(bc_pe_472_io_ve_input),
    .io_input_valid(bc_pe_472_io_input_valid),
    .io_iormac(bc_pe_472_io_iormac),
    .io_ve_out(bc_pe_472_io_ve_out),
    .io_ho_out(bc_pe_472_io_ho_out),
    .io_res_out(bc_pe_472_io_res_out)
  );
  bc_pe bc_pe_473 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_473_clock),
    .reset(bc_pe_473_reset),
    .io_ho_input(bc_pe_473_io_ho_input),
    .io_ve_input(bc_pe_473_io_ve_input),
    .io_input_valid(bc_pe_473_io_input_valid),
    .io_iormac(bc_pe_473_io_iormac),
    .io_ve_out(bc_pe_473_io_ve_out),
    .io_ho_out(bc_pe_473_io_ho_out),
    .io_res_out(bc_pe_473_io_res_out)
  );
  bc_pe bc_pe_474 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_474_clock),
    .reset(bc_pe_474_reset),
    .io_ho_input(bc_pe_474_io_ho_input),
    .io_ve_input(bc_pe_474_io_ve_input),
    .io_input_valid(bc_pe_474_io_input_valid),
    .io_iormac(bc_pe_474_io_iormac),
    .io_ve_out(bc_pe_474_io_ve_out),
    .io_ho_out(bc_pe_474_io_ho_out),
    .io_res_out(bc_pe_474_io_res_out)
  );
  bc_pe bc_pe_475 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_475_clock),
    .reset(bc_pe_475_reset),
    .io_ho_input(bc_pe_475_io_ho_input),
    .io_ve_input(bc_pe_475_io_ve_input),
    .io_input_valid(bc_pe_475_io_input_valid),
    .io_iormac(bc_pe_475_io_iormac),
    .io_ve_out(bc_pe_475_io_ve_out),
    .io_ho_out(bc_pe_475_io_ho_out),
    .io_res_out(bc_pe_475_io_res_out)
  );
  bc_pe bc_pe_476 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_476_clock),
    .reset(bc_pe_476_reset),
    .io_ho_input(bc_pe_476_io_ho_input),
    .io_ve_input(bc_pe_476_io_ve_input),
    .io_input_valid(bc_pe_476_io_input_valid),
    .io_iormac(bc_pe_476_io_iormac),
    .io_ve_out(bc_pe_476_io_ve_out),
    .io_ho_out(bc_pe_476_io_ho_out),
    .io_res_out(bc_pe_476_io_res_out)
  );
  bc_pe bc_pe_477 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_477_clock),
    .reset(bc_pe_477_reset),
    .io_ho_input(bc_pe_477_io_ho_input),
    .io_ve_input(bc_pe_477_io_ve_input),
    .io_input_valid(bc_pe_477_io_input_valid),
    .io_iormac(bc_pe_477_io_iormac),
    .io_ve_out(bc_pe_477_io_ve_out),
    .io_ho_out(bc_pe_477_io_ho_out),
    .io_res_out(bc_pe_477_io_res_out)
  );
  bc_pe bc_pe_478 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_478_clock),
    .reset(bc_pe_478_reset),
    .io_ho_input(bc_pe_478_io_ho_input),
    .io_ve_input(bc_pe_478_io_ve_input),
    .io_input_valid(bc_pe_478_io_input_valid),
    .io_iormac(bc_pe_478_io_iormac),
    .io_ve_out(bc_pe_478_io_ve_out),
    .io_ho_out(bc_pe_478_io_ho_out),
    .io_res_out(bc_pe_478_io_res_out)
  );
  bc_pe bc_pe_479 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_479_clock),
    .reset(bc_pe_479_reset),
    .io_ho_input(bc_pe_479_io_ho_input),
    .io_ve_input(bc_pe_479_io_ve_input),
    .io_input_valid(bc_pe_479_io_input_valid),
    .io_iormac(bc_pe_479_io_iormac),
    .io_ve_out(bc_pe_479_io_ve_out),
    .io_ho_out(bc_pe_479_io_ho_out),
    .io_res_out(bc_pe_479_io_res_out)
  );
  bc_pe bc_pe_480 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_480_clock),
    .reset(bc_pe_480_reset),
    .io_ho_input(bc_pe_480_io_ho_input),
    .io_ve_input(bc_pe_480_io_ve_input),
    .io_input_valid(bc_pe_480_io_input_valid),
    .io_iormac(bc_pe_480_io_iormac),
    .io_ve_out(bc_pe_480_io_ve_out),
    .io_ho_out(bc_pe_480_io_ho_out),
    .io_res_out(bc_pe_480_io_res_out)
  );
  bc_pe bc_pe_481 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_481_clock),
    .reset(bc_pe_481_reset),
    .io_ho_input(bc_pe_481_io_ho_input),
    .io_ve_input(bc_pe_481_io_ve_input),
    .io_input_valid(bc_pe_481_io_input_valid),
    .io_iormac(bc_pe_481_io_iormac),
    .io_ve_out(bc_pe_481_io_ve_out),
    .io_ho_out(bc_pe_481_io_ho_out),
    .io_res_out(bc_pe_481_io_res_out)
  );
  bc_pe bc_pe_482 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_482_clock),
    .reset(bc_pe_482_reset),
    .io_ho_input(bc_pe_482_io_ho_input),
    .io_ve_input(bc_pe_482_io_ve_input),
    .io_input_valid(bc_pe_482_io_input_valid),
    .io_iormac(bc_pe_482_io_iormac),
    .io_ve_out(bc_pe_482_io_ve_out),
    .io_ho_out(bc_pe_482_io_ho_out),
    .io_res_out(bc_pe_482_io_res_out)
  );
  bc_pe bc_pe_483 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_483_clock),
    .reset(bc_pe_483_reset),
    .io_ho_input(bc_pe_483_io_ho_input),
    .io_ve_input(bc_pe_483_io_ve_input),
    .io_input_valid(bc_pe_483_io_input_valid),
    .io_iormac(bc_pe_483_io_iormac),
    .io_ve_out(bc_pe_483_io_ve_out),
    .io_ho_out(bc_pe_483_io_ho_out),
    .io_res_out(bc_pe_483_io_res_out)
  );
  bc_pe bc_pe_484 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_484_clock),
    .reset(bc_pe_484_reset),
    .io_ho_input(bc_pe_484_io_ho_input),
    .io_ve_input(bc_pe_484_io_ve_input),
    .io_input_valid(bc_pe_484_io_input_valid),
    .io_iormac(bc_pe_484_io_iormac),
    .io_ve_out(bc_pe_484_io_ve_out),
    .io_ho_out(bc_pe_484_io_ho_out),
    .io_res_out(bc_pe_484_io_res_out)
  );
  bc_pe bc_pe_485 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_485_clock),
    .reset(bc_pe_485_reset),
    .io_ho_input(bc_pe_485_io_ho_input),
    .io_ve_input(bc_pe_485_io_ve_input),
    .io_input_valid(bc_pe_485_io_input_valid),
    .io_iormac(bc_pe_485_io_iormac),
    .io_ve_out(bc_pe_485_io_ve_out),
    .io_ho_out(bc_pe_485_io_ho_out),
    .io_res_out(bc_pe_485_io_res_out)
  );
  bc_pe bc_pe_486 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_486_clock),
    .reset(bc_pe_486_reset),
    .io_ho_input(bc_pe_486_io_ho_input),
    .io_ve_input(bc_pe_486_io_ve_input),
    .io_input_valid(bc_pe_486_io_input_valid),
    .io_iormac(bc_pe_486_io_iormac),
    .io_ve_out(bc_pe_486_io_ve_out),
    .io_ho_out(bc_pe_486_io_ho_out),
    .io_res_out(bc_pe_486_io_res_out)
  );
  bc_pe bc_pe_487 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_487_clock),
    .reset(bc_pe_487_reset),
    .io_ho_input(bc_pe_487_io_ho_input),
    .io_ve_input(bc_pe_487_io_ve_input),
    .io_input_valid(bc_pe_487_io_input_valid),
    .io_iormac(bc_pe_487_io_iormac),
    .io_ve_out(bc_pe_487_io_ve_out),
    .io_ho_out(bc_pe_487_io_ho_out),
    .io_res_out(bc_pe_487_io_res_out)
  );
  bc_pe bc_pe_488 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_488_clock),
    .reset(bc_pe_488_reset),
    .io_ho_input(bc_pe_488_io_ho_input),
    .io_ve_input(bc_pe_488_io_ve_input),
    .io_input_valid(bc_pe_488_io_input_valid),
    .io_iormac(bc_pe_488_io_iormac),
    .io_ve_out(bc_pe_488_io_ve_out),
    .io_ho_out(bc_pe_488_io_ho_out),
    .io_res_out(bc_pe_488_io_res_out)
  );
  bc_pe bc_pe_489 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_489_clock),
    .reset(bc_pe_489_reset),
    .io_ho_input(bc_pe_489_io_ho_input),
    .io_ve_input(bc_pe_489_io_ve_input),
    .io_input_valid(bc_pe_489_io_input_valid),
    .io_iormac(bc_pe_489_io_iormac),
    .io_ve_out(bc_pe_489_io_ve_out),
    .io_ho_out(bc_pe_489_io_ho_out),
    .io_res_out(bc_pe_489_io_res_out)
  );
  bc_pe bc_pe_490 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_490_clock),
    .reset(bc_pe_490_reset),
    .io_ho_input(bc_pe_490_io_ho_input),
    .io_ve_input(bc_pe_490_io_ve_input),
    .io_input_valid(bc_pe_490_io_input_valid),
    .io_iormac(bc_pe_490_io_iormac),
    .io_ve_out(bc_pe_490_io_ve_out),
    .io_ho_out(bc_pe_490_io_ho_out),
    .io_res_out(bc_pe_490_io_res_out)
  );
  bc_pe bc_pe_491 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_491_clock),
    .reset(bc_pe_491_reset),
    .io_ho_input(bc_pe_491_io_ho_input),
    .io_ve_input(bc_pe_491_io_ve_input),
    .io_input_valid(bc_pe_491_io_input_valid),
    .io_iormac(bc_pe_491_io_iormac),
    .io_ve_out(bc_pe_491_io_ve_out),
    .io_ho_out(bc_pe_491_io_ho_out),
    .io_res_out(bc_pe_491_io_res_out)
  );
  bc_pe bc_pe_492 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_492_clock),
    .reset(bc_pe_492_reset),
    .io_ho_input(bc_pe_492_io_ho_input),
    .io_ve_input(bc_pe_492_io_ve_input),
    .io_input_valid(bc_pe_492_io_input_valid),
    .io_iormac(bc_pe_492_io_iormac),
    .io_ve_out(bc_pe_492_io_ve_out),
    .io_ho_out(bc_pe_492_io_ho_out),
    .io_res_out(bc_pe_492_io_res_out)
  );
  bc_pe bc_pe_493 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_493_clock),
    .reset(bc_pe_493_reset),
    .io_ho_input(bc_pe_493_io_ho_input),
    .io_ve_input(bc_pe_493_io_ve_input),
    .io_input_valid(bc_pe_493_io_input_valid),
    .io_iormac(bc_pe_493_io_iormac),
    .io_ve_out(bc_pe_493_io_ve_out),
    .io_ho_out(bc_pe_493_io_ho_out),
    .io_res_out(bc_pe_493_io_res_out)
  );
  bc_pe bc_pe_494 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_494_clock),
    .reset(bc_pe_494_reset),
    .io_ho_input(bc_pe_494_io_ho_input),
    .io_ve_input(bc_pe_494_io_ve_input),
    .io_input_valid(bc_pe_494_io_input_valid),
    .io_iormac(bc_pe_494_io_iormac),
    .io_ve_out(bc_pe_494_io_ve_out),
    .io_ho_out(bc_pe_494_io_ho_out),
    .io_res_out(bc_pe_494_io_res_out)
  );
  bc_pe bc_pe_495 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_495_clock),
    .reset(bc_pe_495_reset),
    .io_ho_input(bc_pe_495_io_ho_input),
    .io_ve_input(bc_pe_495_io_ve_input),
    .io_input_valid(bc_pe_495_io_input_valid),
    .io_iormac(bc_pe_495_io_iormac),
    .io_ve_out(bc_pe_495_io_ve_out),
    .io_ho_out(bc_pe_495_io_ho_out),
    .io_res_out(bc_pe_495_io_res_out)
  );
  bc_pe bc_pe_496 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_496_clock),
    .reset(bc_pe_496_reset),
    .io_ho_input(bc_pe_496_io_ho_input),
    .io_ve_input(bc_pe_496_io_ve_input),
    .io_input_valid(bc_pe_496_io_input_valid),
    .io_iormac(bc_pe_496_io_iormac),
    .io_ve_out(bc_pe_496_io_ve_out),
    .io_ho_out(bc_pe_496_io_ho_out),
    .io_res_out(bc_pe_496_io_res_out)
  );
  bc_pe bc_pe_497 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_497_clock),
    .reset(bc_pe_497_reset),
    .io_ho_input(bc_pe_497_io_ho_input),
    .io_ve_input(bc_pe_497_io_ve_input),
    .io_input_valid(bc_pe_497_io_input_valid),
    .io_iormac(bc_pe_497_io_iormac),
    .io_ve_out(bc_pe_497_io_ve_out),
    .io_ho_out(bc_pe_497_io_ho_out),
    .io_res_out(bc_pe_497_io_res_out)
  );
  bc_pe bc_pe_498 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_498_clock),
    .reset(bc_pe_498_reset),
    .io_ho_input(bc_pe_498_io_ho_input),
    .io_ve_input(bc_pe_498_io_ve_input),
    .io_input_valid(bc_pe_498_io_input_valid),
    .io_iormac(bc_pe_498_io_iormac),
    .io_ve_out(bc_pe_498_io_ve_out),
    .io_ho_out(bc_pe_498_io_ho_out),
    .io_res_out(bc_pe_498_io_res_out)
  );
  bc_pe bc_pe_499 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_499_clock),
    .reset(bc_pe_499_reset),
    .io_ho_input(bc_pe_499_io_ho_input),
    .io_ve_input(bc_pe_499_io_ve_input),
    .io_input_valid(bc_pe_499_io_input_valid),
    .io_iormac(bc_pe_499_io_iormac),
    .io_ve_out(bc_pe_499_io_ve_out),
    .io_ho_out(bc_pe_499_io_ho_out),
    .io_res_out(bc_pe_499_io_res_out)
  );
  bc_pe bc_pe_500 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_500_clock),
    .reset(bc_pe_500_reset),
    .io_ho_input(bc_pe_500_io_ho_input),
    .io_ve_input(bc_pe_500_io_ve_input),
    .io_input_valid(bc_pe_500_io_input_valid),
    .io_iormac(bc_pe_500_io_iormac),
    .io_ve_out(bc_pe_500_io_ve_out),
    .io_ho_out(bc_pe_500_io_ho_out),
    .io_res_out(bc_pe_500_io_res_out)
  );
  bc_pe bc_pe_501 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_501_clock),
    .reset(bc_pe_501_reset),
    .io_ho_input(bc_pe_501_io_ho_input),
    .io_ve_input(bc_pe_501_io_ve_input),
    .io_input_valid(bc_pe_501_io_input_valid),
    .io_iormac(bc_pe_501_io_iormac),
    .io_ve_out(bc_pe_501_io_ve_out),
    .io_ho_out(bc_pe_501_io_ho_out),
    .io_res_out(bc_pe_501_io_res_out)
  );
  bc_pe bc_pe_502 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_502_clock),
    .reset(bc_pe_502_reset),
    .io_ho_input(bc_pe_502_io_ho_input),
    .io_ve_input(bc_pe_502_io_ve_input),
    .io_input_valid(bc_pe_502_io_input_valid),
    .io_iormac(bc_pe_502_io_iormac),
    .io_ve_out(bc_pe_502_io_ve_out),
    .io_ho_out(bc_pe_502_io_ho_out),
    .io_res_out(bc_pe_502_io_res_out)
  );
  bc_pe bc_pe_503 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_503_clock),
    .reset(bc_pe_503_reset),
    .io_ho_input(bc_pe_503_io_ho_input),
    .io_ve_input(bc_pe_503_io_ve_input),
    .io_input_valid(bc_pe_503_io_input_valid),
    .io_iormac(bc_pe_503_io_iormac),
    .io_ve_out(bc_pe_503_io_ve_out),
    .io_ho_out(bc_pe_503_io_ho_out),
    .io_res_out(bc_pe_503_io_res_out)
  );
  bc_pe bc_pe_504 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_504_clock),
    .reset(bc_pe_504_reset),
    .io_ho_input(bc_pe_504_io_ho_input),
    .io_ve_input(bc_pe_504_io_ve_input),
    .io_input_valid(bc_pe_504_io_input_valid),
    .io_iormac(bc_pe_504_io_iormac),
    .io_ve_out(bc_pe_504_io_ve_out),
    .io_ho_out(bc_pe_504_io_ho_out),
    .io_res_out(bc_pe_504_io_res_out)
  );
  bc_pe bc_pe_505 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_505_clock),
    .reset(bc_pe_505_reset),
    .io_ho_input(bc_pe_505_io_ho_input),
    .io_ve_input(bc_pe_505_io_ve_input),
    .io_input_valid(bc_pe_505_io_input_valid),
    .io_iormac(bc_pe_505_io_iormac),
    .io_ve_out(bc_pe_505_io_ve_out),
    .io_ho_out(bc_pe_505_io_ho_out),
    .io_res_out(bc_pe_505_io_res_out)
  );
  bc_pe bc_pe_506 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_506_clock),
    .reset(bc_pe_506_reset),
    .io_ho_input(bc_pe_506_io_ho_input),
    .io_ve_input(bc_pe_506_io_ve_input),
    .io_input_valid(bc_pe_506_io_input_valid),
    .io_iormac(bc_pe_506_io_iormac),
    .io_ve_out(bc_pe_506_io_ve_out),
    .io_ho_out(bc_pe_506_io_ho_out),
    .io_res_out(bc_pe_506_io_res_out)
  );
  bc_pe bc_pe_507 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_507_clock),
    .reset(bc_pe_507_reset),
    .io_ho_input(bc_pe_507_io_ho_input),
    .io_ve_input(bc_pe_507_io_ve_input),
    .io_input_valid(bc_pe_507_io_input_valid),
    .io_iormac(bc_pe_507_io_iormac),
    .io_ve_out(bc_pe_507_io_ve_out),
    .io_ho_out(bc_pe_507_io_ho_out),
    .io_res_out(bc_pe_507_io_res_out)
  );
  bc_pe bc_pe_508 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_508_clock),
    .reset(bc_pe_508_reset),
    .io_ho_input(bc_pe_508_io_ho_input),
    .io_ve_input(bc_pe_508_io_ve_input),
    .io_input_valid(bc_pe_508_io_input_valid),
    .io_iormac(bc_pe_508_io_iormac),
    .io_ve_out(bc_pe_508_io_ve_out),
    .io_ho_out(bc_pe_508_io_ho_out),
    .io_res_out(bc_pe_508_io_res_out)
  );
  bc_pe bc_pe_509 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_509_clock),
    .reset(bc_pe_509_reset),
    .io_ho_input(bc_pe_509_io_ho_input),
    .io_ve_input(bc_pe_509_io_ve_input),
    .io_input_valid(bc_pe_509_io_input_valid),
    .io_iormac(bc_pe_509_io_iormac),
    .io_ve_out(bc_pe_509_io_ve_out),
    .io_ho_out(bc_pe_509_io_ho_out),
    .io_res_out(bc_pe_509_io_res_out)
  );
  bc_pe bc_pe_510 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_510_clock),
    .reset(bc_pe_510_reset),
    .io_ho_input(bc_pe_510_io_ho_input),
    .io_ve_input(bc_pe_510_io_ve_input),
    .io_input_valid(bc_pe_510_io_input_valid),
    .io_iormac(bc_pe_510_io_iormac),
    .io_ve_out(bc_pe_510_io_ve_out),
    .io_ho_out(bc_pe_510_io_ho_out),
    .io_res_out(bc_pe_510_io_res_out)
  );
  bc_pe bc_pe_511 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_511_clock),
    .reset(bc_pe_511_reset),
    .io_ho_input(bc_pe_511_io_ho_input),
    .io_ve_input(bc_pe_511_io_ve_input),
    .io_input_valid(bc_pe_511_io_input_valid),
    .io_iormac(bc_pe_511_io_iormac),
    .io_ve_out(bc_pe_511_io_ve_out),
    .io_ho_out(bc_pe_511_io_ho_out),
    .io_res_out(bc_pe_511_io_res_out)
  );
  bc_pe bc_pe_512 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_512_clock),
    .reset(bc_pe_512_reset),
    .io_ho_input(bc_pe_512_io_ho_input),
    .io_ve_input(bc_pe_512_io_ve_input),
    .io_input_valid(bc_pe_512_io_input_valid),
    .io_iormac(bc_pe_512_io_iormac),
    .io_ve_out(bc_pe_512_io_ve_out),
    .io_ho_out(bc_pe_512_io_ho_out),
    .io_res_out(bc_pe_512_io_res_out)
  );
  bc_pe bc_pe_513 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_513_clock),
    .reset(bc_pe_513_reset),
    .io_ho_input(bc_pe_513_io_ho_input),
    .io_ve_input(bc_pe_513_io_ve_input),
    .io_input_valid(bc_pe_513_io_input_valid),
    .io_iormac(bc_pe_513_io_iormac),
    .io_ve_out(bc_pe_513_io_ve_out),
    .io_ho_out(bc_pe_513_io_ho_out),
    .io_res_out(bc_pe_513_io_res_out)
  );
  bc_pe bc_pe_514 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_514_clock),
    .reset(bc_pe_514_reset),
    .io_ho_input(bc_pe_514_io_ho_input),
    .io_ve_input(bc_pe_514_io_ve_input),
    .io_input_valid(bc_pe_514_io_input_valid),
    .io_iormac(bc_pe_514_io_iormac),
    .io_ve_out(bc_pe_514_io_ve_out),
    .io_ho_out(bc_pe_514_io_ho_out),
    .io_res_out(bc_pe_514_io_res_out)
  );
  bc_pe bc_pe_515 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_515_clock),
    .reset(bc_pe_515_reset),
    .io_ho_input(bc_pe_515_io_ho_input),
    .io_ve_input(bc_pe_515_io_ve_input),
    .io_input_valid(bc_pe_515_io_input_valid),
    .io_iormac(bc_pe_515_io_iormac),
    .io_ve_out(bc_pe_515_io_ve_out),
    .io_ho_out(bc_pe_515_io_ho_out),
    .io_res_out(bc_pe_515_io_res_out)
  );
  bc_pe bc_pe_516 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_516_clock),
    .reset(bc_pe_516_reset),
    .io_ho_input(bc_pe_516_io_ho_input),
    .io_ve_input(bc_pe_516_io_ve_input),
    .io_input_valid(bc_pe_516_io_input_valid),
    .io_iormac(bc_pe_516_io_iormac),
    .io_ve_out(bc_pe_516_io_ve_out),
    .io_ho_out(bc_pe_516_io_ho_out),
    .io_res_out(bc_pe_516_io_res_out)
  );
  bc_pe bc_pe_517 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_517_clock),
    .reset(bc_pe_517_reset),
    .io_ho_input(bc_pe_517_io_ho_input),
    .io_ve_input(bc_pe_517_io_ve_input),
    .io_input_valid(bc_pe_517_io_input_valid),
    .io_iormac(bc_pe_517_io_iormac),
    .io_ve_out(bc_pe_517_io_ve_out),
    .io_ho_out(bc_pe_517_io_ho_out),
    .io_res_out(bc_pe_517_io_res_out)
  );
  bc_pe bc_pe_518 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_518_clock),
    .reset(bc_pe_518_reset),
    .io_ho_input(bc_pe_518_io_ho_input),
    .io_ve_input(bc_pe_518_io_ve_input),
    .io_input_valid(bc_pe_518_io_input_valid),
    .io_iormac(bc_pe_518_io_iormac),
    .io_ve_out(bc_pe_518_io_ve_out),
    .io_ho_out(bc_pe_518_io_ho_out),
    .io_res_out(bc_pe_518_io_res_out)
  );
  bc_pe bc_pe_519 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_519_clock),
    .reset(bc_pe_519_reset),
    .io_ho_input(bc_pe_519_io_ho_input),
    .io_ve_input(bc_pe_519_io_ve_input),
    .io_input_valid(bc_pe_519_io_input_valid),
    .io_iormac(bc_pe_519_io_iormac),
    .io_ve_out(bc_pe_519_io_ve_out),
    .io_ho_out(bc_pe_519_io_ho_out),
    .io_res_out(bc_pe_519_io_res_out)
  );
  bc_pe bc_pe_520 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_520_clock),
    .reset(bc_pe_520_reset),
    .io_ho_input(bc_pe_520_io_ho_input),
    .io_ve_input(bc_pe_520_io_ve_input),
    .io_input_valid(bc_pe_520_io_input_valid),
    .io_iormac(bc_pe_520_io_iormac),
    .io_ve_out(bc_pe_520_io_ve_out),
    .io_ho_out(bc_pe_520_io_ho_out),
    .io_res_out(bc_pe_520_io_res_out)
  );
  bc_pe bc_pe_521 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_521_clock),
    .reset(bc_pe_521_reset),
    .io_ho_input(bc_pe_521_io_ho_input),
    .io_ve_input(bc_pe_521_io_ve_input),
    .io_input_valid(bc_pe_521_io_input_valid),
    .io_iormac(bc_pe_521_io_iormac),
    .io_ve_out(bc_pe_521_io_ve_out),
    .io_ho_out(bc_pe_521_io_ho_out),
    .io_res_out(bc_pe_521_io_res_out)
  );
  bc_pe bc_pe_522 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_522_clock),
    .reset(bc_pe_522_reset),
    .io_ho_input(bc_pe_522_io_ho_input),
    .io_ve_input(bc_pe_522_io_ve_input),
    .io_input_valid(bc_pe_522_io_input_valid),
    .io_iormac(bc_pe_522_io_iormac),
    .io_ve_out(bc_pe_522_io_ve_out),
    .io_ho_out(bc_pe_522_io_ho_out),
    .io_res_out(bc_pe_522_io_res_out)
  );
  bc_pe bc_pe_523 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_523_clock),
    .reset(bc_pe_523_reset),
    .io_ho_input(bc_pe_523_io_ho_input),
    .io_ve_input(bc_pe_523_io_ve_input),
    .io_input_valid(bc_pe_523_io_input_valid),
    .io_iormac(bc_pe_523_io_iormac),
    .io_ve_out(bc_pe_523_io_ve_out),
    .io_ho_out(bc_pe_523_io_ho_out),
    .io_res_out(bc_pe_523_io_res_out)
  );
  bc_pe bc_pe_524 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_524_clock),
    .reset(bc_pe_524_reset),
    .io_ho_input(bc_pe_524_io_ho_input),
    .io_ve_input(bc_pe_524_io_ve_input),
    .io_input_valid(bc_pe_524_io_input_valid),
    .io_iormac(bc_pe_524_io_iormac),
    .io_ve_out(bc_pe_524_io_ve_out),
    .io_ho_out(bc_pe_524_io_ho_out),
    .io_res_out(bc_pe_524_io_res_out)
  );
  bc_pe bc_pe_525 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_525_clock),
    .reset(bc_pe_525_reset),
    .io_ho_input(bc_pe_525_io_ho_input),
    .io_ve_input(bc_pe_525_io_ve_input),
    .io_input_valid(bc_pe_525_io_input_valid),
    .io_iormac(bc_pe_525_io_iormac),
    .io_ve_out(bc_pe_525_io_ve_out),
    .io_ho_out(bc_pe_525_io_ho_out),
    .io_res_out(bc_pe_525_io_res_out)
  );
  bc_pe bc_pe_526 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_526_clock),
    .reset(bc_pe_526_reset),
    .io_ho_input(bc_pe_526_io_ho_input),
    .io_ve_input(bc_pe_526_io_ve_input),
    .io_input_valid(bc_pe_526_io_input_valid),
    .io_iormac(bc_pe_526_io_iormac),
    .io_ve_out(bc_pe_526_io_ve_out),
    .io_ho_out(bc_pe_526_io_ho_out),
    .io_res_out(bc_pe_526_io_res_out)
  );
  bc_pe bc_pe_527 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_527_clock),
    .reset(bc_pe_527_reset),
    .io_ho_input(bc_pe_527_io_ho_input),
    .io_ve_input(bc_pe_527_io_ve_input),
    .io_input_valid(bc_pe_527_io_input_valid),
    .io_iormac(bc_pe_527_io_iormac),
    .io_ve_out(bc_pe_527_io_ve_out),
    .io_ho_out(bc_pe_527_io_ho_out),
    .io_res_out(bc_pe_527_io_res_out)
  );
  bc_pe bc_pe_528 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_528_clock),
    .reset(bc_pe_528_reset),
    .io_ho_input(bc_pe_528_io_ho_input),
    .io_ve_input(bc_pe_528_io_ve_input),
    .io_input_valid(bc_pe_528_io_input_valid),
    .io_iormac(bc_pe_528_io_iormac),
    .io_ve_out(bc_pe_528_io_ve_out),
    .io_ho_out(bc_pe_528_io_ho_out),
    .io_res_out(bc_pe_528_io_res_out)
  );
  bc_pe bc_pe_529 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_529_clock),
    .reset(bc_pe_529_reset),
    .io_ho_input(bc_pe_529_io_ho_input),
    .io_ve_input(bc_pe_529_io_ve_input),
    .io_input_valid(bc_pe_529_io_input_valid),
    .io_iormac(bc_pe_529_io_iormac),
    .io_ve_out(bc_pe_529_io_ve_out),
    .io_ho_out(bc_pe_529_io_ho_out),
    .io_res_out(bc_pe_529_io_res_out)
  );
  bc_pe bc_pe_530 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_530_clock),
    .reset(bc_pe_530_reset),
    .io_ho_input(bc_pe_530_io_ho_input),
    .io_ve_input(bc_pe_530_io_ve_input),
    .io_input_valid(bc_pe_530_io_input_valid),
    .io_iormac(bc_pe_530_io_iormac),
    .io_ve_out(bc_pe_530_io_ve_out),
    .io_ho_out(bc_pe_530_io_ho_out),
    .io_res_out(bc_pe_530_io_res_out)
  );
  bc_pe bc_pe_531 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_531_clock),
    .reset(bc_pe_531_reset),
    .io_ho_input(bc_pe_531_io_ho_input),
    .io_ve_input(bc_pe_531_io_ve_input),
    .io_input_valid(bc_pe_531_io_input_valid),
    .io_iormac(bc_pe_531_io_iormac),
    .io_ve_out(bc_pe_531_io_ve_out),
    .io_ho_out(bc_pe_531_io_ho_out),
    .io_res_out(bc_pe_531_io_res_out)
  );
  bc_pe bc_pe_532 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_532_clock),
    .reset(bc_pe_532_reset),
    .io_ho_input(bc_pe_532_io_ho_input),
    .io_ve_input(bc_pe_532_io_ve_input),
    .io_input_valid(bc_pe_532_io_input_valid),
    .io_iormac(bc_pe_532_io_iormac),
    .io_ve_out(bc_pe_532_io_ve_out),
    .io_ho_out(bc_pe_532_io_ho_out),
    .io_res_out(bc_pe_532_io_res_out)
  );
  bc_pe bc_pe_533 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_533_clock),
    .reset(bc_pe_533_reset),
    .io_ho_input(bc_pe_533_io_ho_input),
    .io_ve_input(bc_pe_533_io_ve_input),
    .io_input_valid(bc_pe_533_io_input_valid),
    .io_iormac(bc_pe_533_io_iormac),
    .io_ve_out(bc_pe_533_io_ve_out),
    .io_ho_out(bc_pe_533_io_ho_out),
    .io_res_out(bc_pe_533_io_res_out)
  );
  bc_pe bc_pe_534 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_534_clock),
    .reset(bc_pe_534_reset),
    .io_ho_input(bc_pe_534_io_ho_input),
    .io_ve_input(bc_pe_534_io_ve_input),
    .io_input_valid(bc_pe_534_io_input_valid),
    .io_iormac(bc_pe_534_io_iormac),
    .io_ve_out(bc_pe_534_io_ve_out),
    .io_ho_out(bc_pe_534_io_ho_out),
    .io_res_out(bc_pe_534_io_res_out)
  );
  bc_pe bc_pe_535 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_535_clock),
    .reset(bc_pe_535_reset),
    .io_ho_input(bc_pe_535_io_ho_input),
    .io_ve_input(bc_pe_535_io_ve_input),
    .io_input_valid(bc_pe_535_io_input_valid),
    .io_iormac(bc_pe_535_io_iormac),
    .io_ve_out(bc_pe_535_io_ve_out),
    .io_ho_out(bc_pe_535_io_ho_out),
    .io_res_out(bc_pe_535_io_res_out)
  );
  bc_pe bc_pe_536 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_536_clock),
    .reset(bc_pe_536_reset),
    .io_ho_input(bc_pe_536_io_ho_input),
    .io_ve_input(bc_pe_536_io_ve_input),
    .io_input_valid(bc_pe_536_io_input_valid),
    .io_iormac(bc_pe_536_io_iormac),
    .io_ve_out(bc_pe_536_io_ve_out),
    .io_ho_out(bc_pe_536_io_ho_out),
    .io_res_out(bc_pe_536_io_res_out)
  );
  bc_pe bc_pe_537 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_537_clock),
    .reset(bc_pe_537_reset),
    .io_ho_input(bc_pe_537_io_ho_input),
    .io_ve_input(bc_pe_537_io_ve_input),
    .io_input_valid(bc_pe_537_io_input_valid),
    .io_iormac(bc_pe_537_io_iormac),
    .io_ve_out(bc_pe_537_io_ve_out),
    .io_ho_out(bc_pe_537_io_ho_out),
    .io_res_out(bc_pe_537_io_res_out)
  );
  bc_pe bc_pe_538 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_538_clock),
    .reset(bc_pe_538_reset),
    .io_ho_input(bc_pe_538_io_ho_input),
    .io_ve_input(bc_pe_538_io_ve_input),
    .io_input_valid(bc_pe_538_io_input_valid),
    .io_iormac(bc_pe_538_io_iormac),
    .io_ve_out(bc_pe_538_io_ve_out),
    .io_ho_out(bc_pe_538_io_ho_out),
    .io_res_out(bc_pe_538_io_res_out)
  );
  bc_pe bc_pe_539 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_539_clock),
    .reset(bc_pe_539_reset),
    .io_ho_input(bc_pe_539_io_ho_input),
    .io_ve_input(bc_pe_539_io_ve_input),
    .io_input_valid(bc_pe_539_io_input_valid),
    .io_iormac(bc_pe_539_io_iormac),
    .io_ve_out(bc_pe_539_io_ve_out),
    .io_ho_out(bc_pe_539_io_ho_out),
    .io_res_out(bc_pe_539_io_res_out)
  );
  bc_pe bc_pe_540 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_540_clock),
    .reset(bc_pe_540_reset),
    .io_ho_input(bc_pe_540_io_ho_input),
    .io_ve_input(bc_pe_540_io_ve_input),
    .io_input_valid(bc_pe_540_io_input_valid),
    .io_iormac(bc_pe_540_io_iormac),
    .io_ve_out(bc_pe_540_io_ve_out),
    .io_ho_out(bc_pe_540_io_ho_out),
    .io_res_out(bc_pe_540_io_res_out)
  );
  bc_pe bc_pe_541 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_541_clock),
    .reset(bc_pe_541_reset),
    .io_ho_input(bc_pe_541_io_ho_input),
    .io_ve_input(bc_pe_541_io_ve_input),
    .io_input_valid(bc_pe_541_io_input_valid),
    .io_iormac(bc_pe_541_io_iormac),
    .io_ve_out(bc_pe_541_io_ve_out),
    .io_ho_out(bc_pe_541_io_ho_out),
    .io_res_out(bc_pe_541_io_res_out)
  );
  bc_pe bc_pe_542 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_542_clock),
    .reset(bc_pe_542_reset),
    .io_ho_input(bc_pe_542_io_ho_input),
    .io_ve_input(bc_pe_542_io_ve_input),
    .io_input_valid(bc_pe_542_io_input_valid),
    .io_iormac(bc_pe_542_io_iormac),
    .io_ve_out(bc_pe_542_io_ve_out),
    .io_ho_out(bc_pe_542_io_ho_out),
    .io_res_out(bc_pe_542_io_res_out)
  );
  bc_pe bc_pe_543 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_543_clock),
    .reset(bc_pe_543_reset),
    .io_ho_input(bc_pe_543_io_ho_input),
    .io_ve_input(bc_pe_543_io_ve_input),
    .io_input_valid(bc_pe_543_io_input_valid),
    .io_iormac(bc_pe_543_io_iormac),
    .io_ve_out(bc_pe_543_io_ve_out),
    .io_ho_out(bc_pe_543_io_ho_out),
    .io_res_out(bc_pe_543_io_res_out)
  );
  bc_pe bc_pe_544 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_544_clock),
    .reset(bc_pe_544_reset),
    .io_ho_input(bc_pe_544_io_ho_input),
    .io_ve_input(bc_pe_544_io_ve_input),
    .io_input_valid(bc_pe_544_io_input_valid),
    .io_iormac(bc_pe_544_io_iormac),
    .io_ve_out(bc_pe_544_io_ve_out),
    .io_ho_out(bc_pe_544_io_ho_out),
    .io_res_out(bc_pe_544_io_res_out)
  );
  bc_pe bc_pe_545 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_545_clock),
    .reset(bc_pe_545_reset),
    .io_ho_input(bc_pe_545_io_ho_input),
    .io_ve_input(bc_pe_545_io_ve_input),
    .io_input_valid(bc_pe_545_io_input_valid),
    .io_iormac(bc_pe_545_io_iormac),
    .io_ve_out(bc_pe_545_io_ve_out),
    .io_ho_out(bc_pe_545_io_ho_out),
    .io_res_out(bc_pe_545_io_res_out)
  );
  bc_pe bc_pe_546 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_546_clock),
    .reset(bc_pe_546_reset),
    .io_ho_input(bc_pe_546_io_ho_input),
    .io_ve_input(bc_pe_546_io_ve_input),
    .io_input_valid(bc_pe_546_io_input_valid),
    .io_iormac(bc_pe_546_io_iormac),
    .io_ve_out(bc_pe_546_io_ve_out),
    .io_ho_out(bc_pe_546_io_ho_out),
    .io_res_out(bc_pe_546_io_res_out)
  );
  bc_pe bc_pe_547 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_547_clock),
    .reset(bc_pe_547_reset),
    .io_ho_input(bc_pe_547_io_ho_input),
    .io_ve_input(bc_pe_547_io_ve_input),
    .io_input_valid(bc_pe_547_io_input_valid),
    .io_iormac(bc_pe_547_io_iormac),
    .io_ve_out(bc_pe_547_io_ve_out),
    .io_ho_out(bc_pe_547_io_ho_out),
    .io_res_out(bc_pe_547_io_res_out)
  );
  bc_pe bc_pe_548 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_548_clock),
    .reset(bc_pe_548_reset),
    .io_ho_input(bc_pe_548_io_ho_input),
    .io_ve_input(bc_pe_548_io_ve_input),
    .io_input_valid(bc_pe_548_io_input_valid),
    .io_iormac(bc_pe_548_io_iormac),
    .io_ve_out(bc_pe_548_io_ve_out),
    .io_ho_out(bc_pe_548_io_ho_out),
    .io_res_out(bc_pe_548_io_res_out)
  );
  bc_pe bc_pe_549 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_549_clock),
    .reset(bc_pe_549_reset),
    .io_ho_input(bc_pe_549_io_ho_input),
    .io_ve_input(bc_pe_549_io_ve_input),
    .io_input_valid(bc_pe_549_io_input_valid),
    .io_iormac(bc_pe_549_io_iormac),
    .io_ve_out(bc_pe_549_io_ve_out),
    .io_ho_out(bc_pe_549_io_ho_out),
    .io_res_out(bc_pe_549_io_res_out)
  );
  bc_pe bc_pe_550 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_550_clock),
    .reset(bc_pe_550_reset),
    .io_ho_input(bc_pe_550_io_ho_input),
    .io_ve_input(bc_pe_550_io_ve_input),
    .io_input_valid(bc_pe_550_io_input_valid),
    .io_iormac(bc_pe_550_io_iormac),
    .io_ve_out(bc_pe_550_io_ve_out),
    .io_ho_out(bc_pe_550_io_ho_out),
    .io_res_out(bc_pe_550_io_res_out)
  );
  bc_pe bc_pe_551 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_551_clock),
    .reset(bc_pe_551_reset),
    .io_ho_input(bc_pe_551_io_ho_input),
    .io_ve_input(bc_pe_551_io_ve_input),
    .io_input_valid(bc_pe_551_io_input_valid),
    .io_iormac(bc_pe_551_io_iormac),
    .io_ve_out(bc_pe_551_io_ve_out),
    .io_ho_out(bc_pe_551_io_ho_out),
    .io_res_out(bc_pe_551_io_res_out)
  );
  bc_pe bc_pe_552 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_552_clock),
    .reset(bc_pe_552_reset),
    .io_ho_input(bc_pe_552_io_ho_input),
    .io_ve_input(bc_pe_552_io_ve_input),
    .io_input_valid(bc_pe_552_io_input_valid),
    .io_iormac(bc_pe_552_io_iormac),
    .io_ve_out(bc_pe_552_io_ve_out),
    .io_ho_out(bc_pe_552_io_ho_out),
    .io_res_out(bc_pe_552_io_res_out)
  );
  bc_pe bc_pe_553 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_553_clock),
    .reset(bc_pe_553_reset),
    .io_ho_input(bc_pe_553_io_ho_input),
    .io_ve_input(bc_pe_553_io_ve_input),
    .io_input_valid(bc_pe_553_io_input_valid),
    .io_iormac(bc_pe_553_io_iormac),
    .io_ve_out(bc_pe_553_io_ve_out),
    .io_ho_out(bc_pe_553_io_ho_out),
    .io_res_out(bc_pe_553_io_res_out)
  );
  bc_pe bc_pe_554 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_554_clock),
    .reset(bc_pe_554_reset),
    .io_ho_input(bc_pe_554_io_ho_input),
    .io_ve_input(bc_pe_554_io_ve_input),
    .io_input_valid(bc_pe_554_io_input_valid),
    .io_iormac(bc_pe_554_io_iormac),
    .io_ve_out(bc_pe_554_io_ve_out),
    .io_ho_out(bc_pe_554_io_ho_out),
    .io_res_out(bc_pe_554_io_res_out)
  );
  bc_pe bc_pe_555 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_555_clock),
    .reset(bc_pe_555_reset),
    .io_ho_input(bc_pe_555_io_ho_input),
    .io_ve_input(bc_pe_555_io_ve_input),
    .io_input_valid(bc_pe_555_io_input_valid),
    .io_iormac(bc_pe_555_io_iormac),
    .io_ve_out(bc_pe_555_io_ve_out),
    .io_ho_out(bc_pe_555_io_ho_out),
    .io_res_out(bc_pe_555_io_res_out)
  );
  bc_pe bc_pe_556 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_556_clock),
    .reset(bc_pe_556_reset),
    .io_ho_input(bc_pe_556_io_ho_input),
    .io_ve_input(bc_pe_556_io_ve_input),
    .io_input_valid(bc_pe_556_io_input_valid),
    .io_iormac(bc_pe_556_io_iormac),
    .io_ve_out(bc_pe_556_io_ve_out),
    .io_ho_out(bc_pe_556_io_ho_out),
    .io_res_out(bc_pe_556_io_res_out)
  );
  bc_pe bc_pe_557 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_557_clock),
    .reset(bc_pe_557_reset),
    .io_ho_input(bc_pe_557_io_ho_input),
    .io_ve_input(bc_pe_557_io_ve_input),
    .io_input_valid(bc_pe_557_io_input_valid),
    .io_iormac(bc_pe_557_io_iormac),
    .io_ve_out(bc_pe_557_io_ve_out),
    .io_ho_out(bc_pe_557_io_ho_out),
    .io_res_out(bc_pe_557_io_res_out)
  );
  bc_pe bc_pe_558 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_558_clock),
    .reset(bc_pe_558_reset),
    .io_ho_input(bc_pe_558_io_ho_input),
    .io_ve_input(bc_pe_558_io_ve_input),
    .io_input_valid(bc_pe_558_io_input_valid),
    .io_iormac(bc_pe_558_io_iormac),
    .io_ve_out(bc_pe_558_io_ve_out),
    .io_ho_out(bc_pe_558_io_ho_out),
    .io_res_out(bc_pe_558_io_res_out)
  );
  bc_pe bc_pe_559 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_559_clock),
    .reset(bc_pe_559_reset),
    .io_ho_input(bc_pe_559_io_ho_input),
    .io_ve_input(bc_pe_559_io_ve_input),
    .io_input_valid(bc_pe_559_io_input_valid),
    .io_iormac(bc_pe_559_io_iormac),
    .io_ve_out(bc_pe_559_io_ve_out),
    .io_ho_out(bc_pe_559_io_ho_out),
    .io_res_out(bc_pe_559_io_res_out)
  );
  bc_pe bc_pe_560 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_560_clock),
    .reset(bc_pe_560_reset),
    .io_ho_input(bc_pe_560_io_ho_input),
    .io_ve_input(bc_pe_560_io_ve_input),
    .io_input_valid(bc_pe_560_io_input_valid),
    .io_iormac(bc_pe_560_io_iormac),
    .io_ve_out(bc_pe_560_io_ve_out),
    .io_ho_out(bc_pe_560_io_ho_out),
    .io_res_out(bc_pe_560_io_res_out)
  );
  bc_pe bc_pe_561 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_561_clock),
    .reset(bc_pe_561_reset),
    .io_ho_input(bc_pe_561_io_ho_input),
    .io_ve_input(bc_pe_561_io_ve_input),
    .io_input_valid(bc_pe_561_io_input_valid),
    .io_iormac(bc_pe_561_io_iormac),
    .io_ve_out(bc_pe_561_io_ve_out),
    .io_ho_out(bc_pe_561_io_ho_out),
    .io_res_out(bc_pe_561_io_res_out)
  );
  bc_pe bc_pe_562 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_562_clock),
    .reset(bc_pe_562_reset),
    .io_ho_input(bc_pe_562_io_ho_input),
    .io_ve_input(bc_pe_562_io_ve_input),
    .io_input_valid(bc_pe_562_io_input_valid),
    .io_iormac(bc_pe_562_io_iormac),
    .io_ve_out(bc_pe_562_io_ve_out),
    .io_ho_out(bc_pe_562_io_ho_out),
    .io_res_out(bc_pe_562_io_res_out)
  );
  bc_pe bc_pe_563 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_563_clock),
    .reset(bc_pe_563_reset),
    .io_ho_input(bc_pe_563_io_ho_input),
    .io_ve_input(bc_pe_563_io_ve_input),
    .io_input_valid(bc_pe_563_io_input_valid),
    .io_iormac(bc_pe_563_io_iormac),
    .io_ve_out(bc_pe_563_io_ve_out),
    .io_ho_out(bc_pe_563_io_ho_out),
    .io_res_out(bc_pe_563_io_res_out)
  );
  bc_pe bc_pe_564 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_564_clock),
    .reset(bc_pe_564_reset),
    .io_ho_input(bc_pe_564_io_ho_input),
    .io_ve_input(bc_pe_564_io_ve_input),
    .io_input_valid(bc_pe_564_io_input_valid),
    .io_iormac(bc_pe_564_io_iormac),
    .io_ve_out(bc_pe_564_io_ve_out),
    .io_ho_out(bc_pe_564_io_ho_out),
    .io_res_out(bc_pe_564_io_res_out)
  );
  bc_pe bc_pe_565 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_565_clock),
    .reset(bc_pe_565_reset),
    .io_ho_input(bc_pe_565_io_ho_input),
    .io_ve_input(bc_pe_565_io_ve_input),
    .io_input_valid(bc_pe_565_io_input_valid),
    .io_iormac(bc_pe_565_io_iormac),
    .io_ve_out(bc_pe_565_io_ve_out),
    .io_ho_out(bc_pe_565_io_ho_out),
    .io_res_out(bc_pe_565_io_res_out)
  );
  bc_pe bc_pe_566 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_566_clock),
    .reset(bc_pe_566_reset),
    .io_ho_input(bc_pe_566_io_ho_input),
    .io_ve_input(bc_pe_566_io_ve_input),
    .io_input_valid(bc_pe_566_io_input_valid),
    .io_iormac(bc_pe_566_io_iormac),
    .io_ve_out(bc_pe_566_io_ve_out),
    .io_ho_out(bc_pe_566_io_ho_out),
    .io_res_out(bc_pe_566_io_res_out)
  );
  bc_pe bc_pe_567 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_567_clock),
    .reset(bc_pe_567_reset),
    .io_ho_input(bc_pe_567_io_ho_input),
    .io_ve_input(bc_pe_567_io_ve_input),
    .io_input_valid(bc_pe_567_io_input_valid),
    .io_iormac(bc_pe_567_io_iormac),
    .io_ve_out(bc_pe_567_io_ve_out),
    .io_ho_out(bc_pe_567_io_ho_out),
    .io_res_out(bc_pe_567_io_res_out)
  );
  bc_pe bc_pe_568 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_568_clock),
    .reset(bc_pe_568_reset),
    .io_ho_input(bc_pe_568_io_ho_input),
    .io_ve_input(bc_pe_568_io_ve_input),
    .io_input_valid(bc_pe_568_io_input_valid),
    .io_iormac(bc_pe_568_io_iormac),
    .io_ve_out(bc_pe_568_io_ve_out),
    .io_ho_out(bc_pe_568_io_ho_out),
    .io_res_out(bc_pe_568_io_res_out)
  );
  bc_pe bc_pe_569 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_569_clock),
    .reset(bc_pe_569_reset),
    .io_ho_input(bc_pe_569_io_ho_input),
    .io_ve_input(bc_pe_569_io_ve_input),
    .io_input_valid(bc_pe_569_io_input_valid),
    .io_iormac(bc_pe_569_io_iormac),
    .io_ve_out(bc_pe_569_io_ve_out),
    .io_ho_out(bc_pe_569_io_ho_out),
    .io_res_out(bc_pe_569_io_res_out)
  );
  bc_pe bc_pe_570 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_570_clock),
    .reset(bc_pe_570_reset),
    .io_ho_input(bc_pe_570_io_ho_input),
    .io_ve_input(bc_pe_570_io_ve_input),
    .io_input_valid(bc_pe_570_io_input_valid),
    .io_iormac(bc_pe_570_io_iormac),
    .io_ve_out(bc_pe_570_io_ve_out),
    .io_ho_out(bc_pe_570_io_ho_out),
    .io_res_out(bc_pe_570_io_res_out)
  );
  bc_pe bc_pe_571 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_571_clock),
    .reset(bc_pe_571_reset),
    .io_ho_input(bc_pe_571_io_ho_input),
    .io_ve_input(bc_pe_571_io_ve_input),
    .io_input_valid(bc_pe_571_io_input_valid),
    .io_iormac(bc_pe_571_io_iormac),
    .io_ve_out(bc_pe_571_io_ve_out),
    .io_ho_out(bc_pe_571_io_ho_out),
    .io_res_out(bc_pe_571_io_res_out)
  );
  bc_pe bc_pe_572 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_572_clock),
    .reset(bc_pe_572_reset),
    .io_ho_input(bc_pe_572_io_ho_input),
    .io_ve_input(bc_pe_572_io_ve_input),
    .io_input_valid(bc_pe_572_io_input_valid),
    .io_iormac(bc_pe_572_io_iormac),
    .io_ve_out(bc_pe_572_io_ve_out),
    .io_ho_out(bc_pe_572_io_ho_out),
    .io_res_out(bc_pe_572_io_res_out)
  );
  bc_pe bc_pe_573 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_573_clock),
    .reset(bc_pe_573_reset),
    .io_ho_input(bc_pe_573_io_ho_input),
    .io_ve_input(bc_pe_573_io_ve_input),
    .io_input_valid(bc_pe_573_io_input_valid),
    .io_iormac(bc_pe_573_io_iormac),
    .io_ve_out(bc_pe_573_io_ve_out),
    .io_ho_out(bc_pe_573_io_ho_out),
    .io_res_out(bc_pe_573_io_res_out)
  );
  bc_pe bc_pe_574 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_574_clock),
    .reset(bc_pe_574_reset),
    .io_ho_input(bc_pe_574_io_ho_input),
    .io_ve_input(bc_pe_574_io_ve_input),
    .io_input_valid(bc_pe_574_io_input_valid),
    .io_iormac(bc_pe_574_io_iormac),
    .io_ve_out(bc_pe_574_io_ve_out),
    .io_ho_out(bc_pe_574_io_ho_out),
    .io_res_out(bc_pe_574_io_res_out)
  );
  bc_pe bc_pe_575 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_575_clock),
    .reset(bc_pe_575_reset),
    .io_ho_input(bc_pe_575_io_ho_input),
    .io_ve_input(bc_pe_575_io_ve_input),
    .io_input_valid(bc_pe_575_io_input_valid),
    .io_iormac(bc_pe_575_io_iormac),
    .io_ve_out(bc_pe_575_io_ve_out),
    .io_ho_out(bc_pe_575_io_ho_out),
    .io_res_out(bc_pe_575_io_res_out)
  );
  bc_pe bc_pe_576 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_576_clock),
    .reset(bc_pe_576_reset),
    .io_ho_input(bc_pe_576_io_ho_input),
    .io_ve_input(bc_pe_576_io_ve_input),
    .io_input_valid(bc_pe_576_io_input_valid),
    .io_iormac(bc_pe_576_io_iormac),
    .io_ve_out(bc_pe_576_io_ve_out),
    .io_ho_out(bc_pe_576_io_ho_out),
    .io_res_out(bc_pe_576_io_res_out)
  );
  bc_pe bc_pe_577 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_577_clock),
    .reset(bc_pe_577_reset),
    .io_ho_input(bc_pe_577_io_ho_input),
    .io_ve_input(bc_pe_577_io_ve_input),
    .io_input_valid(bc_pe_577_io_input_valid),
    .io_iormac(bc_pe_577_io_iormac),
    .io_ve_out(bc_pe_577_io_ve_out),
    .io_ho_out(bc_pe_577_io_ho_out),
    .io_res_out(bc_pe_577_io_res_out)
  );
  bc_pe bc_pe_578 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_578_clock),
    .reset(bc_pe_578_reset),
    .io_ho_input(bc_pe_578_io_ho_input),
    .io_ve_input(bc_pe_578_io_ve_input),
    .io_input_valid(bc_pe_578_io_input_valid),
    .io_iormac(bc_pe_578_io_iormac),
    .io_ve_out(bc_pe_578_io_ve_out),
    .io_ho_out(bc_pe_578_io_ho_out),
    .io_res_out(bc_pe_578_io_res_out)
  );
  bc_pe bc_pe_579 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_579_clock),
    .reset(bc_pe_579_reset),
    .io_ho_input(bc_pe_579_io_ho_input),
    .io_ve_input(bc_pe_579_io_ve_input),
    .io_input_valid(bc_pe_579_io_input_valid),
    .io_iormac(bc_pe_579_io_iormac),
    .io_ve_out(bc_pe_579_io_ve_out),
    .io_ho_out(bc_pe_579_io_ho_out),
    .io_res_out(bc_pe_579_io_res_out)
  );
  bc_pe bc_pe_580 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_580_clock),
    .reset(bc_pe_580_reset),
    .io_ho_input(bc_pe_580_io_ho_input),
    .io_ve_input(bc_pe_580_io_ve_input),
    .io_input_valid(bc_pe_580_io_input_valid),
    .io_iormac(bc_pe_580_io_iormac),
    .io_ve_out(bc_pe_580_io_ve_out),
    .io_ho_out(bc_pe_580_io_ho_out),
    .io_res_out(bc_pe_580_io_res_out)
  );
  bc_pe bc_pe_581 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_581_clock),
    .reset(bc_pe_581_reset),
    .io_ho_input(bc_pe_581_io_ho_input),
    .io_ve_input(bc_pe_581_io_ve_input),
    .io_input_valid(bc_pe_581_io_input_valid),
    .io_iormac(bc_pe_581_io_iormac),
    .io_ve_out(bc_pe_581_io_ve_out),
    .io_ho_out(bc_pe_581_io_ho_out),
    .io_res_out(bc_pe_581_io_res_out)
  );
  bc_pe bc_pe_582 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_582_clock),
    .reset(bc_pe_582_reset),
    .io_ho_input(bc_pe_582_io_ho_input),
    .io_ve_input(bc_pe_582_io_ve_input),
    .io_input_valid(bc_pe_582_io_input_valid),
    .io_iormac(bc_pe_582_io_iormac),
    .io_ve_out(bc_pe_582_io_ve_out),
    .io_ho_out(bc_pe_582_io_ho_out),
    .io_res_out(bc_pe_582_io_res_out)
  );
  bc_pe bc_pe_583 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_583_clock),
    .reset(bc_pe_583_reset),
    .io_ho_input(bc_pe_583_io_ho_input),
    .io_ve_input(bc_pe_583_io_ve_input),
    .io_input_valid(bc_pe_583_io_input_valid),
    .io_iormac(bc_pe_583_io_iormac),
    .io_ve_out(bc_pe_583_io_ve_out),
    .io_ho_out(bc_pe_583_io_ho_out),
    .io_res_out(bc_pe_583_io_res_out)
  );
  bc_pe bc_pe_584 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_584_clock),
    .reset(bc_pe_584_reset),
    .io_ho_input(bc_pe_584_io_ho_input),
    .io_ve_input(bc_pe_584_io_ve_input),
    .io_input_valid(bc_pe_584_io_input_valid),
    .io_iormac(bc_pe_584_io_iormac),
    .io_ve_out(bc_pe_584_io_ve_out),
    .io_ho_out(bc_pe_584_io_ho_out),
    .io_res_out(bc_pe_584_io_res_out)
  );
  bc_pe bc_pe_585 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_585_clock),
    .reset(bc_pe_585_reset),
    .io_ho_input(bc_pe_585_io_ho_input),
    .io_ve_input(bc_pe_585_io_ve_input),
    .io_input_valid(bc_pe_585_io_input_valid),
    .io_iormac(bc_pe_585_io_iormac),
    .io_ve_out(bc_pe_585_io_ve_out),
    .io_ho_out(bc_pe_585_io_ho_out),
    .io_res_out(bc_pe_585_io_res_out)
  );
  bc_pe bc_pe_586 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_586_clock),
    .reset(bc_pe_586_reset),
    .io_ho_input(bc_pe_586_io_ho_input),
    .io_ve_input(bc_pe_586_io_ve_input),
    .io_input_valid(bc_pe_586_io_input_valid),
    .io_iormac(bc_pe_586_io_iormac),
    .io_ve_out(bc_pe_586_io_ve_out),
    .io_ho_out(bc_pe_586_io_ho_out),
    .io_res_out(bc_pe_586_io_res_out)
  );
  bc_pe bc_pe_587 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_587_clock),
    .reset(bc_pe_587_reset),
    .io_ho_input(bc_pe_587_io_ho_input),
    .io_ve_input(bc_pe_587_io_ve_input),
    .io_input_valid(bc_pe_587_io_input_valid),
    .io_iormac(bc_pe_587_io_iormac),
    .io_ve_out(bc_pe_587_io_ve_out),
    .io_ho_out(bc_pe_587_io_ho_out),
    .io_res_out(bc_pe_587_io_res_out)
  );
  bc_pe bc_pe_588 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_588_clock),
    .reset(bc_pe_588_reset),
    .io_ho_input(bc_pe_588_io_ho_input),
    .io_ve_input(bc_pe_588_io_ve_input),
    .io_input_valid(bc_pe_588_io_input_valid),
    .io_iormac(bc_pe_588_io_iormac),
    .io_ve_out(bc_pe_588_io_ve_out),
    .io_ho_out(bc_pe_588_io_ho_out),
    .io_res_out(bc_pe_588_io_res_out)
  );
  bc_pe bc_pe_589 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_589_clock),
    .reset(bc_pe_589_reset),
    .io_ho_input(bc_pe_589_io_ho_input),
    .io_ve_input(bc_pe_589_io_ve_input),
    .io_input_valid(bc_pe_589_io_input_valid),
    .io_iormac(bc_pe_589_io_iormac),
    .io_ve_out(bc_pe_589_io_ve_out),
    .io_ho_out(bc_pe_589_io_ho_out),
    .io_res_out(bc_pe_589_io_res_out)
  );
  bc_pe bc_pe_590 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_590_clock),
    .reset(bc_pe_590_reset),
    .io_ho_input(bc_pe_590_io_ho_input),
    .io_ve_input(bc_pe_590_io_ve_input),
    .io_input_valid(bc_pe_590_io_input_valid),
    .io_iormac(bc_pe_590_io_iormac),
    .io_ve_out(bc_pe_590_io_ve_out),
    .io_ho_out(bc_pe_590_io_ho_out),
    .io_res_out(bc_pe_590_io_res_out)
  );
  bc_pe bc_pe_591 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_591_clock),
    .reset(bc_pe_591_reset),
    .io_ho_input(bc_pe_591_io_ho_input),
    .io_ve_input(bc_pe_591_io_ve_input),
    .io_input_valid(bc_pe_591_io_input_valid),
    .io_iormac(bc_pe_591_io_iormac),
    .io_ve_out(bc_pe_591_io_ve_out),
    .io_ho_out(bc_pe_591_io_ho_out),
    .io_res_out(bc_pe_591_io_res_out)
  );
  bc_pe bc_pe_592 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_592_clock),
    .reset(bc_pe_592_reset),
    .io_ho_input(bc_pe_592_io_ho_input),
    .io_ve_input(bc_pe_592_io_ve_input),
    .io_input_valid(bc_pe_592_io_input_valid),
    .io_iormac(bc_pe_592_io_iormac),
    .io_ve_out(bc_pe_592_io_ve_out),
    .io_ho_out(bc_pe_592_io_ho_out),
    .io_res_out(bc_pe_592_io_res_out)
  );
  bc_pe bc_pe_593 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_593_clock),
    .reset(bc_pe_593_reset),
    .io_ho_input(bc_pe_593_io_ho_input),
    .io_ve_input(bc_pe_593_io_ve_input),
    .io_input_valid(bc_pe_593_io_input_valid),
    .io_iormac(bc_pe_593_io_iormac),
    .io_ve_out(bc_pe_593_io_ve_out),
    .io_ho_out(bc_pe_593_io_ho_out),
    .io_res_out(bc_pe_593_io_res_out)
  );
  bc_pe bc_pe_594 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_594_clock),
    .reset(bc_pe_594_reset),
    .io_ho_input(bc_pe_594_io_ho_input),
    .io_ve_input(bc_pe_594_io_ve_input),
    .io_input_valid(bc_pe_594_io_input_valid),
    .io_iormac(bc_pe_594_io_iormac),
    .io_ve_out(bc_pe_594_io_ve_out),
    .io_ho_out(bc_pe_594_io_ho_out),
    .io_res_out(bc_pe_594_io_res_out)
  );
  bc_pe bc_pe_595 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_595_clock),
    .reset(bc_pe_595_reset),
    .io_ho_input(bc_pe_595_io_ho_input),
    .io_ve_input(bc_pe_595_io_ve_input),
    .io_input_valid(bc_pe_595_io_input_valid),
    .io_iormac(bc_pe_595_io_iormac),
    .io_ve_out(bc_pe_595_io_ve_out),
    .io_ho_out(bc_pe_595_io_ho_out),
    .io_res_out(bc_pe_595_io_res_out)
  );
  bc_pe bc_pe_596 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_596_clock),
    .reset(bc_pe_596_reset),
    .io_ho_input(bc_pe_596_io_ho_input),
    .io_ve_input(bc_pe_596_io_ve_input),
    .io_input_valid(bc_pe_596_io_input_valid),
    .io_iormac(bc_pe_596_io_iormac),
    .io_ve_out(bc_pe_596_io_ve_out),
    .io_ho_out(bc_pe_596_io_ho_out),
    .io_res_out(bc_pe_596_io_res_out)
  );
  bc_pe bc_pe_597 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_597_clock),
    .reset(bc_pe_597_reset),
    .io_ho_input(bc_pe_597_io_ho_input),
    .io_ve_input(bc_pe_597_io_ve_input),
    .io_input_valid(bc_pe_597_io_input_valid),
    .io_iormac(bc_pe_597_io_iormac),
    .io_ve_out(bc_pe_597_io_ve_out),
    .io_ho_out(bc_pe_597_io_ho_out),
    .io_res_out(bc_pe_597_io_res_out)
  );
  bc_pe bc_pe_598 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_598_clock),
    .reset(bc_pe_598_reset),
    .io_ho_input(bc_pe_598_io_ho_input),
    .io_ve_input(bc_pe_598_io_ve_input),
    .io_input_valid(bc_pe_598_io_input_valid),
    .io_iormac(bc_pe_598_io_iormac),
    .io_ve_out(bc_pe_598_io_ve_out),
    .io_ho_out(bc_pe_598_io_ho_out),
    .io_res_out(bc_pe_598_io_res_out)
  );
  bc_pe bc_pe_599 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_599_clock),
    .reset(bc_pe_599_reset),
    .io_ho_input(bc_pe_599_io_ho_input),
    .io_ve_input(bc_pe_599_io_ve_input),
    .io_input_valid(bc_pe_599_io_input_valid),
    .io_iormac(bc_pe_599_io_iormac),
    .io_ve_out(bc_pe_599_io_ve_out),
    .io_ho_out(bc_pe_599_io_ho_out),
    .io_res_out(bc_pe_599_io_res_out)
  );
  bc_pe bc_pe_600 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_600_clock),
    .reset(bc_pe_600_reset),
    .io_ho_input(bc_pe_600_io_ho_input),
    .io_ve_input(bc_pe_600_io_ve_input),
    .io_input_valid(bc_pe_600_io_input_valid),
    .io_iormac(bc_pe_600_io_iormac),
    .io_ve_out(bc_pe_600_io_ve_out),
    .io_ho_out(bc_pe_600_io_ho_out),
    .io_res_out(bc_pe_600_io_res_out)
  );
  bc_pe bc_pe_601 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_601_clock),
    .reset(bc_pe_601_reset),
    .io_ho_input(bc_pe_601_io_ho_input),
    .io_ve_input(bc_pe_601_io_ve_input),
    .io_input_valid(bc_pe_601_io_input_valid),
    .io_iormac(bc_pe_601_io_iormac),
    .io_ve_out(bc_pe_601_io_ve_out),
    .io_ho_out(bc_pe_601_io_ho_out),
    .io_res_out(bc_pe_601_io_res_out)
  );
  bc_pe bc_pe_602 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_602_clock),
    .reset(bc_pe_602_reset),
    .io_ho_input(bc_pe_602_io_ho_input),
    .io_ve_input(bc_pe_602_io_ve_input),
    .io_input_valid(bc_pe_602_io_input_valid),
    .io_iormac(bc_pe_602_io_iormac),
    .io_ve_out(bc_pe_602_io_ve_out),
    .io_ho_out(bc_pe_602_io_ho_out),
    .io_res_out(bc_pe_602_io_res_out)
  );
  bc_pe bc_pe_603 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_603_clock),
    .reset(bc_pe_603_reset),
    .io_ho_input(bc_pe_603_io_ho_input),
    .io_ve_input(bc_pe_603_io_ve_input),
    .io_input_valid(bc_pe_603_io_input_valid),
    .io_iormac(bc_pe_603_io_iormac),
    .io_ve_out(bc_pe_603_io_ve_out),
    .io_ho_out(bc_pe_603_io_ho_out),
    .io_res_out(bc_pe_603_io_res_out)
  );
  bc_pe bc_pe_604 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_604_clock),
    .reset(bc_pe_604_reset),
    .io_ho_input(bc_pe_604_io_ho_input),
    .io_ve_input(bc_pe_604_io_ve_input),
    .io_input_valid(bc_pe_604_io_input_valid),
    .io_iormac(bc_pe_604_io_iormac),
    .io_ve_out(bc_pe_604_io_ve_out),
    .io_ho_out(bc_pe_604_io_ho_out),
    .io_res_out(bc_pe_604_io_res_out)
  );
  bc_pe bc_pe_605 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_605_clock),
    .reset(bc_pe_605_reset),
    .io_ho_input(bc_pe_605_io_ho_input),
    .io_ve_input(bc_pe_605_io_ve_input),
    .io_input_valid(bc_pe_605_io_input_valid),
    .io_iormac(bc_pe_605_io_iormac),
    .io_ve_out(bc_pe_605_io_ve_out),
    .io_ho_out(bc_pe_605_io_ho_out),
    .io_res_out(bc_pe_605_io_res_out)
  );
  bc_pe bc_pe_606 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_606_clock),
    .reset(bc_pe_606_reset),
    .io_ho_input(bc_pe_606_io_ho_input),
    .io_ve_input(bc_pe_606_io_ve_input),
    .io_input_valid(bc_pe_606_io_input_valid),
    .io_iormac(bc_pe_606_io_iormac),
    .io_ve_out(bc_pe_606_io_ve_out),
    .io_ho_out(bc_pe_606_io_ho_out),
    .io_res_out(bc_pe_606_io_res_out)
  );
  bc_pe bc_pe_607 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_607_clock),
    .reset(bc_pe_607_reset),
    .io_ho_input(bc_pe_607_io_ho_input),
    .io_ve_input(bc_pe_607_io_ve_input),
    .io_input_valid(bc_pe_607_io_input_valid),
    .io_iormac(bc_pe_607_io_iormac),
    .io_ve_out(bc_pe_607_io_ve_out),
    .io_ho_out(bc_pe_607_io_ho_out),
    .io_res_out(bc_pe_607_io_res_out)
  );
  bc_pe bc_pe_608 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_608_clock),
    .reset(bc_pe_608_reset),
    .io_ho_input(bc_pe_608_io_ho_input),
    .io_ve_input(bc_pe_608_io_ve_input),
    .io_input_valid(bc_pe_608_io_input_valid),
    .io_iormac(bc_pe_608_io_iormac),
    .io_ve_out(bc_pe_608_io_ve_out),
    .io_ho_out(bc_pe_608_io_ho_out),
    .io_res_out(bc_pe_608_io_res_out)
  );
  bc_pe bc_pe_609 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_609_clock),
    .reset(bc_pe_609_reset),
    .io_ho_input(bc_pe_609_io_ho_input),
    .io_ve_input(bc_pe_609_io_ve_input),
    .io_input_valid(bc_pe_609_io_input_valid),
    .io_iormac(bc_pe_609_io_iormac),
    .io_ve_out(bc_pe_609_io_ve_out),
    .io_ho_out(bc_pe_609_io_ho_out),
    .io_res_out(bc_pe_609_io_res_out)
  );
  bc_pe bc_pe_610 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_610_clock),
    .reset(bc_pe_610_reset),
    .io_ho_input(bc_pe_610_io_ho_input),
    .io_ve_input(bc_pe_610_io_ve_input),
    .io_input_valid(bc_pe_610_io_input_valid),
    .io_iormac(bc_pe_610_io_iormac),
    .io_ve_out(bc_pe_610_io_ve_out),
    .io_ho_out(bc_pe_610_io_ho_out),
    .io_res_out(bc_pe_610_io_res_out)
  );
  bc_pe bc_pe_611 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_611_clock),
    .reset(bc_pe_611_reset),
    .io_ho_input(bc_pe_611_io_ho_input),
    .io_ve_input(bc_pe_611_io_ve_input),
    .io_input_valid(bc_pe_611_io_input_valid),
    .io_iormac(bc_pe_611_io_iormac),
    .io_ve_out(bc_pe_611_io_ve_out),
    .io_ho_out(bc_pe_611_io_ho_out),
    .io_res_out(bc_pe_611_io_res_out)
  );
  bc_pe bc_pe_612 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_612_clock),
    .reset(bc_pe_612_reset),
    .io_ho_input(bc_pe_612_io_ho_input),
    .io_ve_input(bc_pe_612_io_ve_input),
    .io_input_valid(bc_pe_612_io_input_valid),
    .io_iormac(bc_pe_612_io_iormac),
    .io_ve_out(bc_pe_612_io_ve_out),
    .io_ho_out(bc_pe_612_io_ho_out),
    .io_res_out(bc_pe_612_io_res_out)
  );
  bc_pe bc_pe_613 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_613_clock),
    .reset(bc_pe_613_reset),
    .io_ho_input(bc_pe_613_io_ho_input),
    .io_ve_input(bc_pe_613_io_ve_input),
    .io_input_valid(bc_pe_613_io_input_valid),
    .io_iormac(bc_pe_613_io_iormac),
    .io_ve_out(bc_pe_613_io_ve_out),
    .io_ho_out(bc_pe_613_io_ho_out),
    .io_res_out(bc_pe_613_io_res_out)
  );
  bc_pe bc_pe_614 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_614_clock),
    .reset(bc_pe_614_reset),
    .io_ho_input(bc_pe_614_io_ho_input),
    .io_ve_input(bc_pe_614_io_ve_input),
    .io_input_valid(bc_pe_614_io_input_valid),
    .io_iormac(bc_pe_614_io_iormac),
    .io_ve_out(bc_pe_614_io_ve_out),
    .io_ho_out(bc_pe_614_io_ho_out),
    .io_res_out(bc_pe_614_io_res_out)
  );
  bc_pe bc_pe_615 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_615_clock),
    .reset(bc_pe_615_reset),
    .io_ho_input(bc_pe_615_io_ho_input),
    .io_ve_input(bc_pe_615_io_ve_input),
    .io_input_valid(bc_pe_615_io_input_valid),
    .io_iormac(bc_pe_615_io_iormac),
    .io_ve_out(bc_pe_615_io_ve_out),
    .io_ho_out(bc_pe_615_io_ho_out),
    .io_res_out(bc_pe_615_io_res_out)
  );
  bc_pe bc_pe_616 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_616_clock),
    .reset(bc_pe_616_reset),
    .io_ho_input(bc_pe_616_io_ho_input),
    .io_ve_input(bc_pe_616_io_ve_input),
    .io_input_valid(bc_pe_616_io_input_valid),
    .io_iormac(bc_pe_616_io_iormac),
    .io_ve_out(bc_pe_616_io_ve_out),
    .io_ho_out(bc_pe_616_io_ho_out),
    .io_res_out(bc_pe_616_io_res_out)
  );
  bc_pe bc_pe_617 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_617_clock),
    .reset(bc_pe_617_reset),
    .io_ho_input(bc_pe_617_io_ho_input),
    .io_ve_input(bc_pe_617_io_ve_input),
    .io_input_valid(bc_pe_617_io_input_valid),
    .io_iormac(bc_pe_617_io_iormac),
    .io_ve_out(bc_pe_617_io_ve_out),
    .io_ho_out(bc_pe_617_io_ho_out),
    .io_res_out(bc_pe_617_io_res_out)
  );
  bc_pe bc_pe_618 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_618_clock),
    .reset(bc_pe_618_reset),
    .io_ho_input(bc_pe_618_io_ho_input),
    .io_ve_input(bc_pe_618_io_ve_input),
    .io_input_valid(bc_pe_618_io_input_valid),
    .io_iormac(bc_pe_618_io_iormac),
    .io_ve_out(bc_pe_618_io_ve_out),
    .io_ho_out(bc_pe_618_io_ho_out),
    .io_res_out(bc_pe_618_io_res_out)
  );
  bc_pe bc_pe_619 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_619_clock),
    .reset(bc_pe_619_reset),
    .io_ho_input(bc_pe_619_io_ho_input),
    .io_ve_input(bc_pe_619_io_ve_input),
    .io_input_valid(bc_pe_619_io_input_valid),
    .io_iormac(bc_pe_619_io_iormac),
    .io_ve_out(bc_pe_619_io_ve_out),
    .io_ho_out(bc_pe_619_io_ho_out),
    .io_res_out(bc_pe_619_io_res_out)
  );
  bc_pe bc_pe_620 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_620_clock),
    .reset(bc_pe_620_reset),
    .io_ho_input(bc_pe_620_io_ho_input),
    .io_ve_input(bc_pe_620_io_ve_input),
    .io_input_valid(bc_pe_620_io_input_valid),
    .io_iormac(bc_pe_620_io_iormac),
    .io_ve_out(bc_pe_620_io_ve_out),
    .io_ho_out(bc_pe_620_io_ho_out),
    .io_res_out(bc_pe_620_io_res_out)
  );
  bc_pe bc_pe_621 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_621_clock),
    .reset(bc_pe_621_reset),
    .io_ho_input(bc_pe_621_io_ho_input),
    .io_ve_input(bc_pe_621_io_ve_input),
    .io_input_valid(bc_pe_621_io_input_valid),
    .io_iormac(bc_pe_621_io_iormac),
    .io_ve_out(bc_pe_621_io_ve_out),
    .io_ho_out(bc_pe_621_io_ho_out),
    .io_res_out(bc_pe_621_io_res_out)
  );
  bc_pe bc_pe_622 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_622_clock),
    .reset(bc_pe_622_reset),
    .io_ho_input(bc_pe_622_io_ho_input),
    .io_ve_input(bc_pe_622_io_ve_input),
    .io_input_valid(bc_pe_622_io_input_valid),
    .io_iormac(bc_pe_622_io_iormac),
    .io_ve_out(bc_pe_622_io_ve_out),
    .io_ho_out(bc_pe_622_io_ho_out),
    .io_res_out(bc_pe_622_io_res_out)
  );
  bc_pe bc_pe_623 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_623_clock),
    .reset(bc_pe_623_reset),
    .io_ho_input(bc_pe_623_io_ho_input),
    .io_ve_input(bc_pe_623_io_ve_input),
    .io_input_valid(bc_pe_623_io_input_valid),
    .io_iormac(bc_pe_623_io_iormac),
    .io_ve_out(bc_pe_623_io_ve_out),
    .io_ho_out(bc_pe_623_io_ho_out),
    .io_res_out(bc_pe_623_io_res_out)
  );
  bc_pe bc_pe_624 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_624_clock),
    .reset(bc_pe_624_reset),
    .io_ho_input(bc_pe_624_io_ho_input),
    .io_ve_input(bc_pe_624_io_ve_input),
    .io_input_valid(bc_pe_624_io_input_valid),
    .io_iormac(bc_pe_624_io_iormac),
    .io_ve_out(bc_pe_624_io_ve_out),
    .io_ho_out(bc_pe_624_io_ho_out),
    .io_res_out(bc_pe_624_io_res_out)
  );
  bc_pe bc_pe_625 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_625_clock),
    .reset(bc_pe_625_reset),
    .io_ho_input(bc_pe_625_io_ho_input),
    .io_ve_input(bc_pe_625_io_ve_input),
    .io_input_valid(bc_pe_625_io_input_valid),
    .io_iormac(bc_pe_625_io_iormac),
    .io_ve_out(bc_pe_625_io_ve_out),
    .io_ho_out(bc_pe_625_io_ho_out),
    .io_res_out(bc_pe_625_io_res_out)
  );
  bc_pe bc_pe_626 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_626_clock),
    .reset(bc_pe_626_reset),
    .io_ho_input(bc_pe_626_io_ho_input),
    .io_ve_input(bc_pe_626_io_ve_input),
    .io_input_valid(bc_pe_626_io_input_valid),
    .io_iormac(bc_pe_626_io_iormac),
    .io_ve_out(bc_pe_626_io_ve_out),
    .io_ho_out(bc_pe_626_io_ho_out),
    .io_res_out(bc_pe_626_io_res_out)
  );
  bc_pe bc_pe_627 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_627_clock),
    .reset(bc_pe_627_reset),
    .io_ho_input(bc_pe_627_io_ho_input),
    .io_ve_input(bc_pe_627_io_ve_input),
    .io_input_valid(bc_pe_627_io_input_valid),
    .io_iormac(bc_pe_627_io_iormac),
    .io_ve_out(bc_pe_627_io_ve_out),
    .io_ho_out(bc_pe_627_io_ho_out),
    .io_res_out(bc_pe_627_io_res_out)
  );
  bc_pe bc_pe_628 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_628_clock),
    .reset(bc_pe_628_reset),
    .io_ho_input(bc_pe_628_io_ho_input),
    .io_ve_input(bc_pe_628_io_ve_input),
    .io_input_valid(bc_pe_628_io_input_valid),
    .io_iormac(bc_pe_628_io_iormac),
    .io_ve_out(bc_pe_628_io_ve_out),
    .io_ho_out(bc_pe_628_io_ho_out),
    .io_res_out(bc_pe_628_io_res_out)
  );
  bc_pe bc_pe_629 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_629_clock),
    .reset(bc_pe_629_reset),
    .io_ho_input(bc_pe_629_io_ho_input),
    .io_ve_input(bc_pe_629_io_ve_input),
    .io_input_valid(bc_pe_629_io_input_valid),
    .io_iormac(bc_pe_629_io_iormac),
    .io_ve_out(bc_pe_629_io_ve_out),
    .io_ho_out(bc_pe_629_io_ho_out),
    .io_res_out(bc_pe_629_io_res_out)
  );
  bc_pe bc_pe_630 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_630_clock),
    .reset(bc_pe_630_reset),
    .io_ho_input(bc_pe_630_io_ho_input),
    .io_ve_input(bc_pe_630_io_ve_input),
    .io_input_valid(bc_pe_630_io_input_valid),
    .io_iormac(bc_pe_630_io_iormac),
    .io_ve_out(bc_pe_630_io_ve_out),
    .io_ho_out(bc_pe_630_io_ho_out),
    .io_res_out(bc_pe_630_io_res_out)
  );
  bc_pe bc_pe_631 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_631_clock),
    .reset(bc_pe_631_reset),
    .io_ho_input(bc_pe_631_io_ho_input),
    .io_ve_input(bc_pe_631_io_ve_input),
    .io_input_valid(bc_pe_631_io_input_valid),
    .io_iormac(bc_pe_631_io_iormac),
    .io_ve_out(bc_pe_631_io_ve_out),
    .io_ho_out(bc_pe_631_io_ho_out),
    .io_res_out(bc_pe_631_io_res_out)
  );
  bc_pe bc_pe_632 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_632_clock),
    .reset(bc_pe_632_reset),
    .io_ho_input(bc_pe_632_io_ho_input),
    .io_ve_input(bc_pe_632_io_ve_input),
    .io_input_valid(bc_pe_632_io_input_valid),
    .io_iormac(bc_pe_632_io_iormac),
    .io_ve_out(bc_pe_632_io_ve_out),
    .io_ho_out(bc_pe_632_io_ho_out),
    .io_res_out(bc_pe_632_io_res_out)
  );
  bc_pe bc_pe_633 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_633_clock),
    .reset(bc_pe_633_reset),
    .io_ho_input(bc_pe_633_io_ho_input),
    .io_ve_input(bc_pe_633_io_ve_input),
    .io_input_valid(bc_pe_633_io_input_valid),
    .io_iormac(bc_pe_633_io_iormac),
    .io_ve_out(bc_pe_633_io_ve_out),
    .io_ho_out(bc_pe_633_io_ho_out),
    .io_res_out(bc_pe_633_io_res_out)
  );
  bc_pe bc_pe_634 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_634_clock),
    .reset(bc_pe_634_reset),
    .io_ho_input(bc_pe_634_io_ho_input),
    .io_ve_input(bc_pe_634_io_ve_input),
    .io_input_valid(bc_pe_634_io_input_valid),
    .io_iormac(bc_pe_634_io_iormac),
    .io_ve_out(bc_pe_634_io_ve_out),
    .io_ho_out(bc_pe_634_io_ho_out),
    .io_res_out(bc_pe_634_io_res_out)
  );
  bc_pe bc_pe_635 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_635_clock),
    .reset(bc_pe_635_reset),
    .io_ho_input(bc_pe_635_io_ho_input),
    .io_ve_input(bc_pe_635_io_ve_input),
    .io_input_valid(bc_pe_635_io_input_valid),
    .io_iormac(bc_pe_635_io_iormac),
    .io_ve_out(bc_pe_635_io_ve_out),
    .io_ho_out(bc_pe_635_io_ho_out),
    .io_res_out(bc_pe_635_io_res_out)
  );
  bc_pe bc_pe_636 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_636_clock),
    .reset(bc_pe_636_reset),
    .io_ho_input(bc_pe_636_io_ho_input),
    .io_ve_input(bc_pe_636_io_ve_input),
    .io_input_valid(bc_pe_636_io_input_valid),
    .io_iormac(bc_pe_636_io_iormac),
    .io_ve_out(bc_pe_636_io_ve_out),
    .io_ho_out(bc_pe_636_io_ho_out),
    .io_res_out(bc_pe_636_io_res_out)
  );
  bc_pe bc_pe_637 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_637_clock),
    .reset(bc_pe_637_reset),
    .io_ho_input(bc_pe_637_io_ho_input),
    .io_ve_input(bc_pe_637_io_ve_input),
    .io_input_valid(bc_pe_637_io_input_valid),
    .io_iormac(bc_pe_637_io_iormac),
    .io_ve_out(bc_pe_637_io_ve_out),
    .io_ho_out(bc_pe_637_io_ho_out),
    .io_res_out(bc_pe_637_io_res_out)
  );
  bc_pe bc_pe_638 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_638_clock),
    .reset(bc_pe_638_reset),
    .io_ho_input(bc_pe_638_io_ho_input),
    .io_ve_input(bc_pe_638_io_ve_input),
    .io_input_valid(bc_pe_638_io_input_valid),
    .io_iormac(bc_pe_638_io_iormac),
    .io_ve_out(bc_pe_638_io_ve_out),
    .io_ho_out(bc_pe_638_io_ho_out),
    .io_res_out(bc_pe_638_io_res_out)
  );
  bc_pe bc_pe_639 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_639_clock),
    .reset(bc_pe_639_reset),
    .io_ho_input(bc_pe_639_io_ho_input),
    .io_ve_input(bc_pe_639_io_ve_input),
    .io_input_valid(bc_pe_639_io_input_valid),
    .io_iormac(bc_pe_639_io_iormac),
    .io_ve_out(bc_pe_639_io_ve_out),
    .io_ho_out(bc_pe_639_io_ho_out),
    .io_res_out(bc_pe_639_io_res_out)
  );
  bc_pe bc_pe_640 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_640_clock),
    .reset(bc_pe_640_reset),
    .io_ho_input(bc_pe_640_io_ho_input),
    .io_ve_input(bc_pe_640_io_ve_input),
    .io_input_valid(bc_pe_640_io_input_valid),
    .io_iormac(bc_pe_640_io_iormac),
    .io_ve_out(bc_pe_640_io_ve_out),
    .io_ho_out(bc_pe_640_io_ho_out),
    .io_res_out(bc_pe_640_io_res_out)
  );
  bc_pe bc_pe_641 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_641_clock),
    .reset(bc_pe_641_reset),
    .io_ho_input(bc_pe_641_io_ho_input),
    .io_ve_input(bc_pe_641_io_ve_input),
    .io_input_valid(bc_pe_641_io_input_valid),
    .io_iormac(bc_pe_641_io_iormac),
    .io_ve_out(bc_pe_641_io_ve_out),
    .io_ho_out(bc_pe_641_io_ho_out),
    .io_res_out(bc_pe_641_io_res_out)
  );
  bc_pe bc_pe_642 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_642_clock),
    .reset(bc_pe_642_reset),
    .io_ho_input(bc_pe_642_io_ho_input),
    .io_ve_input(bc_pe_642_io_ve_input),
    .io_input_valid(bc_pe_642_io_input_valid),
    .io_iormac(bc_pe_642_io_iormac),
    .io_ve_out(bc_pe_642_io_ve_out),
    .io_ho_out(bc_pe_642_io_ho_out),
    .io_res_out(bc_pe_642_io_res_out)
  );
  bc_pe bc_pe_643 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_643_clock),
    .reset(bc_pe_643_reset),
    .io_ho_input(bc_pe_643_io_ho_input),
    .io_ve_input(bc_pe_643_io_ve_input),
    .io_input_valid(bc_pe_643_io_input_valid),
    .io_iormac(bc_pe_643_io_iormac),
    .io_ve_out(bc_pe_643_io_ve_out),
    .io_ho_out(bc_pe_643_io_ho_out),
    .io_res_out(bc_pe_643_io_res_out)
  );
  bc_pe bc_pe_644 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_644_clock),
    .reset(bc_pe_644_reset),
    .io_ho_input(bc_pe_644_io_ho_input),
    .io_ve_input(bc_pe_644_io_ve_input),
    .io_input_valid(bc_pe_644_io_input_valid),
    .io_iormac(bc_pe_644_io_iormac),
    .io_ve_out(bc_pe_644_io_ve_out),
    .io_ho_out(bc_pe_644_io_ho_out),
    .io_res_out(bc_pe_644_io_res_out)
  );
  bc_pe bc_pe_645 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_645_clock),
    .reset(bc_pe_645_reset),
    .io_ho_input(bc_pe_645_io_ho_input),
    .io_ve_input(bc_pe_645_io_ve_input),
    .io_input_valid(bc_pe_645_io_input_valid),
    .io_iormac(bc_pe_645_io_iormac),
    .io_ve_out(bc_pe_645_io_ve_out),
    .io_ho_out(bc_pe_645_io_ho_out),
    .io_res_out(bc_pe_645_io_res_out)
  );
  bc_pe bc_pe_646 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_646_clock),
    .reset(bc_pe_646_reset),
    .io_ho_input(bc_pe_646_io_ho_input),
    .io_ve_input(bc_pe_646_io_ve_input),
    .io_input_valid(bc_pe_646_io_input_valid),
    .io_iormac(bc_pe_646_io_iormac),
    .io_ve_out(bc_pe_646_io_ve_out),
    .io_ho_out(bc_pe_646_io_ho_out),
    .io_res_out(bc_pe_646_io_res_out)
  );
  bc_pe bc_pe_647 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_647_clock),
    .reset(bc_pe_647_reset),
    .io_ho_input(bc_pe_647_io_ho_input),
    .io_ve_input(bc_pe_647_io_ve_input),
    .io_input_valid(bc_pe_647_io_input_valid),
    .io_iormac(bc_pe_647_io_iormac),
    .io_ve_out(bc_pe_647_io_ve_out),
    .io_ho_out(bc_pe_647_io_ho_out),
    .io_res_out(bc_pe_647_io_res_out)
  );
  bc_pe bc_pe_648 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_648_clock),
    .reset(bc_pe_648_reset),
    .io_ho_input(bc_pe_648_io_ho_input),
    .io_ve_input(bc_pe_648_io_ve_input),
    .io_input_valid(bc_pe_648_io_input_valid),
    .io_iormac(bc_pe_648_io_iormac),
    .io_ve_out(bc_pe_648_io_ve_out),
    .io_ho_out(bc_pe_648_io_ho_out),
    .io_res_out(bc_pe_648_io_res_out)
  );
  bc_pe bc_pe_649 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_649_clock),
    .reset(bc_pe_649_reset),
    .io_ho_input(bc_pe_649_io_ho_input),
    .io_ve_input(bc_pe_649_io_ve_input),
    .io_input_valid(bc_pe_649_io_input_valid),
    .io_iormac(bc_pe_649_io_iormac),
    .io_ve_out(bc_pe_649_io_ve_out),
    .io_ho_out(bc_pe_649_io_ho_out),
    .io_res_out(bc_pe_649_io_res_out)
  );
  bc_pe bc_pe_650 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_650_clock),
    .reset(bc_pe_650_reset),
    .io_ho_input(bc_pe_650_io_ho_input),
    .io_ve_input(bc_pe_650_io_ve_input),
    .io_input_valid(bc_pe_650_io_input_valid),
    .io_iormac(bc_pe_650_io_iormac),
    .io_ve_out(bc_pe_650_io_ve_out),
    .io_ho_out(bc_pe_650_io_ho_out),
    .io_res_out(bc_pe_650_io_res_out)
  );
  bc_pe bc_pe_651 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_651_clock),
    .reset(bc_pe_651_reset),
    .io_ho_input(bc_pe_651_io_ho_input),
    .io_ve_input(bc_pe_651_io_ve_input),
    .io_input_valid(bc_pe_651_io_input_valid),
    .io_iormac(bc_pe_651_io_iormac),
    .io_ve_out(bc_pe_651_io_ve_out),
    .io_ho_out(bc_pe_651_io_ho_out),
    .io_res_out(bc_pe_651_io_res_out)
  );
  bc_pe bc_pe_652 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_652_clock),
    .reset(bc_pe_652_reset),
    .io_ho_input(bc_pe_652_io_ho_input),
    .io_ve_input(bc_pe_652_io_ve_input),
    .io_input_valid(bc_pe_652_io_input_valid),
    .io_iormac(bc_pe_652_io_iormac),
    .io_ve_out(bc_pe_652_io_ve_out),
    .io_ho_out(bc_pe_652_io_ho_out),
    .io_res_out(bc_pe_652_io_res_out)
  );
  bc_pe bc_pe_653 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_653_clock),
    .reset(bc_pe_653_reset),
    .io_ho_input(bc_pe_653_io_ho_input),
    .io_ve_input(bc_pe_653_io_ve_input),
    .io_input_valid(bc_pe_653_io_input_valid),
    .io_iormac(bc_pe_653_io_iormac),
    .io_ve_out(bc_pe_653_io_ve_out),
    .io_ho_out(bc_pe_653_io_ho_out),
    .io_res_out(bc_pe_653_io_res_out)
  );
  bc_pe bc_pe_654 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_654_clock),
    .reset(bc_pe_654_reset),
    .io_ho_input(bc_pe_654_io_ho_input),
    .io_ve_input(bc_pe_654_io_ve_input),
    .io_input_valid(bc_pe_654_io_input_valid),
    .io_iormac(bc_pe_654_io_iormac),
    .io_ve_out(bc_pe_654_io_ve_out),
    .io_ho_out(bc_pe_654_io_ho_out),
    .io_res_out(bc_pe_654_io_res_out)
  );
  bc_pe bc_pe_655 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_655_clock),
    .reset(bc_pe_655_reset),
    .io_ho_input(bc_pe_655_io_ho_input),
    .io_ve_input(bc_pe_655_io_ve_input),
    .io_input_valid(bc_pe_655_io_input_valid),
    .io_iormac(bc_pe_655_io_iormac),
    .io_ve_out(bc_pe_655_io_ve_out),
    .io_ho_out(bc_pe_655_io_ho_out),
    .io_res_out(bc_pe_655_io_res_out)
  );
  bc_pe bc_pe_656 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_656_clock),
    .reset(bc_pe_656_reset),
    .io_ho_input(bc_pe_656_io_ho_input),
    .io_ve_input(bc_pe_656_io_ve_input),
    .io_input_valid(bc_pe_656_io_input_valid),
    .io_iormac(bc_pe_656_io_iormac),
    .io_ve_out(bc_pe_656_io_ve_out),
    .io_ho_out(bc_pe_656_io_ho_out),
    .io_res_out(bc_pe_656_io_res_out)
  );
  bc_pe bc_pe_657 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_657_clock),
    .reset(bc_pe_657_reset),
    .io_ho_input(bc_pe_657_io_ho_input),
    .io_ve_input(bc_pe_657_io_ve_input),
    .io_input_valid(bc_pe_657_io_input_valid),
    .io_iormac(bc_pe_657_io_iormac),
    .io_ve_out(bc_pe_657_io_ve_out),
    .io_ho_out(bc_pe_657_io_ho_out),
    .io_res_out(bc_pe_657_io_res_out)
  );
  bc_pe bc_pe_658 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_658_clock),
    .reset(bc_pe_658_reset),
    .io_ho_input(bc_pe_658_io_ho_input),
    .io_ve_input(bc_pe_658_io_ve_input),
    .io_input_valid(bc_pe_658_io_input_valid),
    .io_iormac(bc_pe_658_io_iormac),
    .io_ve_out(bc_pe_658_io_ve_out),
    .io_ho_out(bc_pe_658_io_ho_out),
    .io_res_out(bc_pe_658_io_res_out)
  );
  bc_pe bc_pe_659 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_659_clock),
    .reset(bc_pe_659_reset),
    .io_ho_input(bc_pe_659_io_ho_input),
    .io_ve_input(bc_pe_659_io_ve_input),
    .io_input_valid(bc_pe_659_io_input_valid),
    .io_iormac(bc_pe_659_io_iormac),
    .io_ve_out(bc_pe_659_io_ve_out),
    .io_ho_out(bc_pe_659_io_ho_out),
    .io_res_out(bc_pe_659_io_res_out)
  );
  bc_pe bc_pe_660 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_660_clock),
    .reset(bc_pe_660_reset),
    .io_ho_input(bc_pe_660_io_ho_input),
    .io_ve_input(bc_pe_660_io_ve_input),
    .io_input_valid(bc_pe_660_io_input_valid),
    .io_iormac(bc_pe_660_io_iormac),
    .io_ve_out(bc_pe_660_io_ve_out),
    .io_ho_out(bc_pe_660_io_ho_out),
    .io_res_out(bc_pe_660_io_res_out)
  );
  bc_pe bc_pe_661 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_661_clock),
    .reset(bc_pe_661_reset),
    .io_ho_input(bc_pe_661_io_ho_input),
    .io_ve_input(bc_pe_661_io_ve_input),
    .io_input_valid(bc_pe_661_io_input_valid),
    .io_iormac(bc_pe_661_io_iormac),
    .io_ve_out(bc_pe_661_io_ve_out),
    .io_ho_out(bc_pe_661_io_ho_out),
    .io_res_out(bc_pe_661_io_res_out)
  );
  bc_pe bc_pe_662 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_662_clock),
    .reset(bc_pe_662_reset),
    .io_ho_input(bc_pe_662_io_ho_input),
    .io_ve_input(bc_pe_662_io_ve_input),
    .io_input_valid(bc_pe_662_io_input_valid),
    .io_iormac(bc_pe_662_io_iormac),
    .io_ve_out(bc_pe_662_io_ve_out),
    .io_ho_out(bc_pe_662_io_ho_out),
    .io_res_out(bc_pe_662_io_res_out)
  );
  bc_pe bc_pe_663 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_663_clock),
    .reset(bc_pe_663_reset),
    .io_ho_input(bc_pe_663_io_ho_input),
    .io_ve_input(bc_pe_663_io_ve_input),
    .io_input_valid(bc_pe_663_io_input_valid),
    .io_iormac(bc_pe_663_io_iormac),
    .io_ve_out(bc_pe_663_io_ve_out),
    .io_ho_out(bc_pe_663_io_ho_out),
    .io_res_out(bc_pe_663_io_res_out)
  );
  bc_pe bc_pe_664 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_664_clock),
    .reset(bc_pe_664_reset),
    .io_ho_input(bc_pe_664_io_ho_input),
    .io_ve_input(bc_pe_664_io_ve_input),
    .io_input_valid(bc_pe_664_io_input_valid),
    .io_iormac(bc_pe_664_io_iormac),
    .io_ve_out(bc_pe_664_io_ve_out),
    .io_ho_out(bc_pe_664_io_ho_out),
    .io_res_out(bc_pe_664_io_res_out)
  );
  bc_pe bc_pe_665 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_665_clock),
    .reset(bc_pe_665_reset),
    .io_ho_input(bc_pe_665_io_ho_input),
    .io_ve_input(bc_pe_665_io_ve_input),
    .io_input_valid(bc_pe_665_io_input_valid),
    .io_iormac(bc_pe_665_io_iormac),
    .io_ve_out(bc_pe_665_io_ve_out),
    .io_ho_out(bc_pe_665_io_ho_out),
    .io_res_out(bc_pe_665_io_res_out)
  );
  bc_pe bc_pe_666 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_666_clock),
    .reset(bc_pe_666_reset),
    .io_ho_input(bc_pe_666_io_ho_input),
    .io_ve_input(bc_pe_666_io_ve_input),
    .io_input_valid(bc_pe_666_io_input_valid),
    .io_iormac(bc_pe_666_io_iormac),
    .io_ve_out(bc_pe_666_io_ve_out),
    .io_ho_out(bc_pe_666_io_ho_out),
    .io_res_out(bc_pe_666_io_res_out)
  );
  bc_pe bc_pe_667 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_667_clock),
    .reset(bc_pe_667_reset),
    .io_ho_input(bc_pe_667_io_ho_input),
    .io_ve_input(bc_pe_667_io_ve_input),
    .io_input_valid(bc_pe_667_io_input_valid),
    .io_iormac(bc_pe_667_io_iormac),
    .io_ve_out(bc_pe_667_io_ve_out),
    .io_ho_out(bc_pe_667_io_ho_out),
    .io_res_out(bc_pe_667_io_res_out)
  );
  bc_pe bc_pe_668 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_668_clock),
    .reset(bc_pe_668_reset),
    .io_ho_input(bc_pe_668_io_ho_input),
    .io_ve_input(bc_pe_668_io_ve_input),
    .io_input_valid(bc_pe_668_io_input_valid),
    .io_iormac(bc_pe_668_io_iormac),
    .io_ve_out(bc_pe_668_io_ve_out),
    .io_ho_out(bc_pe_668_io_ho_out),
    .io_res_out(bc_pe_668_io_res_out)
  );
  bc_pe bc_pe_669 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_669_clock),
    .reset(bc_pe_669_reset),
    .io_ho_input(bc_pe_669_io_ho_input),
    .io_ve_input(bc_pe_669_io_ve_input),
    .io_input_valid(bc_pe_669_io_input_valid),
    .io_iormac(bc_pe_669_io_iormac),
    .io_ve_out(bc_pe_669_io_ve_out),
    .io_ho_out(bc_pe_669_io_ho_out),
    .io_res_out(bc_pe_669_io_res_out)
  );
  bc_pe bc_pe_670 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_670_clock),
    .reset(bc_pe_670_reset),
    .io_ho_input(bc_pe_670_io_ho_input),
    .io_ve_input(bc_pe_670_io_ve_input),
    .io_input_valid(bc_pe_670_io_input_valid),
    .io_iormac(bc_pe_670_io_iormac),
    .io_ve_out(bc_pe_670_io_ve_out),
    .io_ho_out(bc_pe_670_io_ho_out),
    .io_res_out(bc_pe_670_io_res_out)
  );
  bc_pe bc_pe_671 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_671_clock),
    .reset(bc_pe_671_reset),
    .io_ho_input(bc_pe_671_io_ho_input),
    .io_ve_input(bc_pe_671_io_ve_input),
    .io_input_valid(bc_pe_671_io_input_valid),
    .io_iormac(bc_pe_671_io_iormac),
    .io_ve_out(bc_pe_671_io_ve_out),
    .io_ho_out(bc_pe_671_io_ho_out),
    .io_res_out(bc_pe_671_io_res_out)
  );
  bc_pe bc_pe_672 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_672_clock),
    .reset(bc_pe_672_reset),
    .io_ho_input(bc_pe_672_io_ho_input),
    .io_ve_input(bc_pe_672_io_ve_input),
    .io_input_valid(bc_pe_672_io_input_valid),
    .io_iormac(bc_pe_672_io_iormac),
    .io_ve_out(bc_pe_672_io_ve_out),
    .io_ho_out(bc_pe_672_io_ho_out),
    .io_res_out(bc_pe_672_io_res_out)
  );
  bc_pe bc_pe_673 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_673_clock),
    .reset(bc_pe_673_reset),
    .io_ho_input(bc_pe_673_io_ho_input),
    .io_ve_input(bc_pe_673_io_ve_input),
    .io_input_valid(bc_pe_673_io_input_valid),
    .io_iormac(bc_pe_673_io_iormac),
    .io_ve_out(bc_pe_673_io_ve_out),
    .io_ho_out(bc_pe_673_io_ho_out),
    .io_res_out(bc_pe_673_io_res_out)
  );
  bc_pe bc_pe_674 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_674_clock),
    .reset(bc_pe_674_reset),
    .io_ho_input(bc_pe_674_io_ho_input),
    .io_ve_input(bc_pe_674_io_ve_input),
    .io_input_valid(bc_pe_674_io_input_valid),
    .io_iormac(bc_pe_674_io_iormac),
    .io_ve_out(bc_pe_674_io_ve_out),
    .io_ho_out(bc_pe_674_io_ho_out),
    .io_res_out(bc_pe_674_io_res_out)
  );
  bc_pe bc_pe_675 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_675_clock),
    .reset(bc_pe_675_reset),
    .io_ho_input(bc_pe_675_io_ho_input),
    .io_ve_input(bc_pe_675_io_ve_input),
    .io_input_valid(bc_pe_675_io_input_valid),
    .io_iormac(bc_pe_675_io_iormac),
    .io_ve_out(bc_pe_675_io_ve_out),
    .io_ho_out(bc_pe_675_io_ho_out),
    .io_res_out(bc_pe_675_io_res_out)
  );
  bc_pe bc_pe_676 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_676_clock),
    .reset(bc_pe_676_reset),
    .io_ho_input(bc_pe_676_io_ho_input),
    .io_ve_input(bc_pe_676_io_ve_input),
    .io_input_valid(bc_pe_676_io_input_valid),
    .io_iormac(bc_pe_676_io_iormac),
    .io_ve_out(bc_pe_676_io_ve_out),
    .io_ho_out(bc_pe_676_io_ho_out),
    .io_res_out(bc_pe_676_io_res_out)
  );
  bc_pe bc_pe_677 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_677_clock),
    .reset(bc_pe_677_reset),
    .io_ho_input(bc_pe_677_io_ho_input),
    .io_ve_input(bc_pe_677_io_ve_input),
    .io_input_valid(bc_pe_677_io_input_valid),
    .io_iormac(bc_pe_677_io_iormac),
    .io_ve_out(bc_pe_677_io_ve_out),
    .io_ho_out(bc_pe_677_io_ho_out),
    .io_res_out(bc_pe_677_io_res_out)
  );
  bc_pe bc_pe_678 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_678_clock),
    .reset(bc_pe_678_reset),
    .io_ho_input(bc_pe_678_io_ho_input),
    .io_ve_input(bc_pe_678_io_ve_input),
    .io_input_valid(bc_pe_678_io_input_valid),
    .io_iormac(bc_pe_678_io_iormac),
    .io_ve_out(bc_pe_678_io_ve_out),
    .io_ho_out(bc_pe_678_io_ho_out),
    .io_res_out(bc_pe_678_io_res_out)
  );
  bc_pe bc_pe_679 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_679_clock),
    .reset(bc_pe_679_reset),
    .io_ho_input(bc_pe_679_io_ho_input),
    .io_ve_input(bc_pe_679_io_ve_input),
    .io_input_valid(bc_pe_679_io_input_valid),
    .io_iormac(bc_pe_679_io_iormac),
    .io_ve_out(bc_pe_679_io_ve_out),
    .io_ho_out(bc_pe_679_io_ho_out),
    .io_res_out(bc_pe_679_io_res_out)
  );
  bc_pe bc_pe_680 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_680_clock),
    .reset(bc_pe_680_reset),
    .io_ho_input(bc_pe_680_io_ho_input),
    .io_ve_input(bc_pe_680_io_ve_input),
    .io_input_valid(bc_pe_680_io_input_valid),
    .io_iormac(bc_pe_680_io_iormac),
    .io_ve_out(bc_pe_680_io_ve_out),
    .io_ho_out(bc_pe_680_io_ho_out),
    .io_res_out(bc_pe_680_io_res_out)
  );
  bc_pe bc_pe_681 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_681_clock),
    .reset(bc_pe_681_reset),
    .io_ho_input(bc_pe_681_io_ho_input),
    .io_ve_input(bc_pe_681_io_ve_input),
    .io_input_valid(bc_pe_681_io_input_valid),
    .io_iormac(bc_pe_681_io_iormac),
    .io_ve_out(bc_pe_681_io_ve_out),
    .io_ho_out(bc_pe_681_io_ho_out),
    .io_res_out(bc_pe_681_io_res_out)
  );
  bc_pe bc_pe_682 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_682_clock),
    .reset(bc_pe_682_reset),
    .io_ho_input(bc_pe_682_io_ho_input),
    .io_ve_input(bc_pe_682_io_ve_input),
    .io_input_valid(bc_pe_682_io_input_valid),
    .io_iormac(bc_pe_682_io_iormac),
    .io_ve_out(bc_pe_682_io_ve_out),
    .io_ho_out(bc_pe_682_io_ho_out),
    .io_res_out(bc_pe_682_io_res_out)
  );
  bc_pe bc_pe_683 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_683_clock),
    .reset(bc_pe_683_reset),
    .io_ho_input(bc_pe_683_io_ho_input),
    .io_ve_input(bc_pe_683_io_ve_input),
    .io_input_valid(bc_pe_683_io_input_valid),
    .io_iormac(bc_pe_683_io_iormac),
    .io_ve_out(bc_pe_683_io_ve_out),
    .io_ho_out(bc_pe_683_io_ho_out),
    .io_res_out(bc_pe_683_io_res_out)
  );
  bc_pe bc_pe_684 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_684_clock),
    .reset(bc_pe_684_reset),
    .io_ho_input(bc_pe_684_io_ho_input),
    .io_ve_input(bc_pe_684_io_ve_input),
    .io_input_valid(bc_pe_684_io_input_valid),
    .io_iormac(bc_pe_684_io_iormac),
    .io_ve_out(bc_pe_684_io_ve_out),
    .io_ho_out(bc_pe_684_io_ho_out),
    .io_res_out(bc_pe_684_io_res_out)
  );
  bc_pe bc_pe_685 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_685_clock),
    .reset(bc_pe_685_reset),
    .io_ho_input(bc_pe_685_io_ho_input),
    .io_ve_input(bc_pe_685_io_ve_input),
    .io_input_valid(bc_pe_685_io_input_valid),
    .io_iormac(bc_pe_685_io_iormac),
    .io_ve_out(bc_pe_685_io_ve_out),
    .io_ho_out(bc_pe_685_io_ho_out),
    .io_res_out(bc_pe_685_io_res_out)
  );
  bc_pe bc_pe_686 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_686_clock),
    .reset(bc_pe_686_reset),
    .io_ho_input(bc_pe_686_io_ho_input),
    .io_ve_input(bc_pe_686_io_ve_input),
    .io_input_valid(bc_pe_686_io_input_valid),
    .io_iormac(bc_pe_686_io_iormac),
    .io_ve_out(bc_pe_686_io_ve_out),
    .io_ho_out(bc_pe_686_io_ho_out),
    .io_res_out(bc_pe_686_io_res_out)
  );
  bc_pe bc_pe_687 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_687_clock),
    .reset(bc_pe_687_reset),
    .io_ho_input(bc_pe_687_io_ho_input),
    .io_ve_input(bc_pe_687_io_ve_input),
    .io_input_valid(bc_pe_687_io_input_valid),
    .io_iormac(bc_pe_687_io_iormac),
    .io_ve_out(bc_pe_687_io_ve_out),
    .io_ho_out(bc_pe_687_io_ho_out),
    .io_res_out(bc_pe_687_io_res_out)
  );
  bc_pe bc_pe_688 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_688_clock),
    .reset(bc_pe_688_reset),
    .io_ho_input(bc_pe_688_io_ho_input),
    .io_ve_input(bc_pe_688_io_ve_input),
    .io_input_valid(bc_pe_688_io_input_valid),
    .io_iormac(bc_pe_688_io_iormac),
    .io_ve_out(bc_pe_688_io_ve_out),
    .io_ho_out(bc_pe_688_io_ho_out),
    .io_res_out(bc_pe_688_io_res_out)
  );
  bc_pe bc_pe_689 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_689_clock),
    .reset(bc_pe_689_reset),
    .io_ho_input(bc_pe_689_io_ho_input),
    .io_ve_input(bc_pe_689_io_ve_input),
    .io_input_valid(bc_pe_689_io_input_valid),
    .io_iormac(bc_pe_689_io_iormac),
    .io_ve_out(bc_pe_689_io_ve_out),
    .io_ho_out(bc_pe_689_io_ho_out),
    .io_res_out(bc_pe_689_io_res_out)
  );
  bc_pe bc_pe_690 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_690_clock),
    .reset(bc_pe_690_reset),
    .io_ho_input(bc_pe_690_io_ho_input),
    .io_ve_input(bc_pe_690_io_ve_input),
    .io_input_valid(bc_pe_690_io_input_valid),
    .io_iormac(bc_pe_690_io_iormac),
    .io_ve_out(bc_pe_690_io_ve_out),
    .io_ho_out(bc_pe_690_io_ho_out),
    .io_res_out(bc_pe_690_io_res_out)
  );
  bc_pe bc_pe_691 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_691_clock),
    .reset(bc_pe_691_reset),
    .io_ho_input(bc_pe_691_io_ho_input),
    .io_ve_input(bc_pe_691_io_ve_input),
    .io_input_valid(bc_pe_691_io_input_valid),
    .io_iormac(bc_pe_691_io_iormac),
    .io_ve_out(bc_pe_691_io_ve_out),
    .io_ho_out(bc_pe_691_io_ho_out),
    .io_res_out(bc_pe_691_io_res_out)
  );
  bc_pe bc_pe_692 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_692_clock),
    .reset(bc_pe_692_reset),
    .io_ho_input(bc_pe_692_io_ho_input),
    .io_ve_input(bc_pe_692_io_ve_input),
    .io_input_valid(bc_pe_692_io_input_valid),
    .io_iormac(bc_pe_692_io_iormac),
    .io_ve_out(bc_pe_692_io_ve_out),
    .io_ho_out(bc_pe_692_io_ho_out),
    .io_res_out(bc_pe_692_io_res_out)
  );
  bc_pe bc_pe_693 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_693_clock),
    .reset(bc_pe_693_reset),
    .io_ho_input(bc_pe_693_io_ho_input),
    .io_ve_input(bc_pe_693_io_ve_input),
    .io_input_valid(bc_pe_693_io_input_valid),
    .io_iormac(bc_pe_693_io_iormac),
    .io_ve_out(bc_pe_693_io_ve_out),
    .io_ho_out(bc_pe_693_io_ho_out),
    .io_res_out(bc_pe_693_io_res_out)
  );
  bc_pe bc_pe_694 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_694_clock),
    .reset(bc_pe_694_reset),
    .io_ho_input(bc_pe_694_io_ho_input),
    .io_ve_input(bc_pe_694_io_ve_input),
    .io_input_valid(bc_pe_694_io_input_valid),
    .io_iormac(bc_pe_694_io_iormac),
    .io_ve_out(bc_pe_694_io_ve_out),
    .io_ho_out(bc_pe_694_io_ho_out),
    .io_res_out(bc_pe_694_io_res_out)
  );
  bc_pe bc_pe_695 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_695_clock),
    .reset(bc_pe_695_reset),
    .io_ho_input(bc_pe_695_io_ho_input),
    .io_ve_input(bc_pe_695_io_ve_input),
    .io_input_valid(bc_pe_695_io_input_valid),
    .io_iormac(bc_pe_695_io_iormac),
    .io_ve_out(bc_pe_695_io_ve_out),
    .io_ho_out(bc_pe_695_io_ho_out),
    .io_res_out(bc_pe_695_io_res_out)
  );
  bc_pe bc_pe_696 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_696_clock),
    .reset(bc_pe_696_reset),
    .io_ho_input(bc_pe_696_io_ho_input),
    .io_ve_input(bc_pe_696_io_ve_input),
    .io_input_valid(bc_pe_696_io_input_valid),
    .io_iormac(bc_pe_696_io_iormac),
    .io_ve_out(bc_pe_696_io_ve_out),
    .io_ho_out(bc_pe_696_io_ho_out),
    .io_res_out(bc_pe_696_io_res_out)
  );
  bc_pe bc_pe_697 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_697_clock),
    .reset(bc_pe_697_reset),
    .io_ho_input(bc_pe_697_io_ho_input),
    .io_ve_input(bc_pe_697_io_ve_input),
    .io_input_valid(bc_pe_697_io_input_valid),
    .io_iormac(bc_pe_697_io_iormac),
    .io_ve_out(bc_pe_697_io_ve_out),
    .io_ho_out(bc_pe_697_io_ho_out),
    .io_res_out(bc_pe_697_io_res_out)
  );
  bc_pe bc_pe_698 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_698_clock),
    .reset(bc_pe_698_reset),
    .io_ho_input(bc_pe_698_io_ho_input),
    .io_ve_input(bc_pe_698_io_ve_input),
    .io_input_valid(bc_pe_698_io_input_valid),
    .io_iormac(bc_pe_698_io_iormac),
    .io_ve_out(bc_pe_698_io_ve_out),
    .io_ho_out(bc_pe_698_io_ho_out),
    .io_res_out(bc_pe_698_io_res_out)
  );
  bc_pe bc_pe_699 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_699_clock),
    .reset(bc_pe_699_reset),
    .io_ho_input(bc_pe_699_io_ho_input),
    .io_ve_input(bc_pe_699_io_ve_input),
    .io_input_valid(bc_pe_699_io_input_valid),
    .io_iormac(bc_pe_699_io_iormac),
    .io_ve_out(bc_pe_699_io_ve_out),
    .io_ho_out(bc_pe_699_io_ho_out),
    .io_res_out(bc_pe_699_io_res_out)
  );
  bc_pe bc_pe_700 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_700_clock),
    .reset(bc_pe_700_reset),
    .io_ho_input(bc_pe_700_io_ho_input),
    .io_ve_input(bc_pe_700_io_ve_input),
    .io_input_valid(bc_pe_700_io_input_valid),
    .io_iormac(bc_pe_700_io_iormac),
    .io_ve_out(bc_pe_700_io_ve_out),
    .io_ho_out(bc_pe_700_io_ho_out),
    .io_res_out(bc_pe_700_io_res_out)
  );
  bc_pe bc_pe_701 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_701_clock),
    .reset(bc_pe_701_reset),
    .io_ho_input(bc_pe_701_io_ho_input),
    .io_ve_input(bc_pe_701_io_ve_input),
    .io_input_valid(bc_pe_701_io_input_valid),
    .io_iormac(bc_pe_701_io_iormac),
    .io_ve_out(bc_pe_701_io_ve_out),
    .io_ho_out(bc_pe_701_io_ho_out),
    .io_res_out(bc_pe_701_io_res_out)
  );
  bc_pe bc_pe_702 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_702_clock),
    .reset(bc_pe_702_reset),
    .io_ho_input(bc_pe_702_io_ho_input),
    .io_ve_input(bc_pe_702_io_ve_input),
    .io_input_valid(bc_pe_702_io_input_valid),
    .io_iormac(bc_pe_702_io_iormac),
    .io_ve_out(bc_pe_702_io_ve_out),
    .io_ho_out(bc_pe_702_io_ho_out),
    .io_res_out(bc_pe_702_io_res_out)
  );
  bc_pe bc_pe_703 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_703_clock),
    .reset(bc_pe_703_reset),
    .io_ho_input(bc_pe_703_io_ho_input),
    .io_ve_input(bc_pe_703_io_ve_input),
    .io_input_valid(bc_pe_703_io_input_valid),
    .io_iormac(bc_pe_703_io_iormac),
    .io_ve_out(bc_pe_703_io_ve_out),
    .io_ho_out(bc_pe_703_io_ho_out),
    .io_res_out(bc_pe_703_io_res_out)
  );
  bc_pe bc_pe_704 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_704_clock),
    .reset(bc_pe_704_reset),
    .io_ho_input(bc_pe_704_io_ho_input),
    .io_ve_input(bc_pe_704_io_ve_input),
    .io_input_valid(bc_pe_704_io_input_valid),
    .io_iormac(bc_pe_704_io_iormac),
    .io_ve_out(bc_pe_704_io_ve_out),
    .io_ho_out(bc_pe_704_io_ho_out),
    .io_res_out(bc_pe_704_io_res_out)
  );
  bc_pe bc_pe_705 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_705_clock),
    .reset(bc_pe_705_reset),
    .io_ho_input(bc_pe_705_io_ho_input),
    .io_ve_input(bc_pe_705_io_ve_input),
    .io_input_valid(bc_pe_705_io_input_valid),
    .io_iormac(bc_pe_705_io_iormac),
    .io_ve_out(bc_pe_705_io_ve_out),
    .io_ho_out(bc_pe_705_io_ho_out),
    .io_res_out(bc_pe_705_io_res_out)
  );
  bc_pe bc_pe_706 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_706_clock),
    .reset(bc_pe_706_reset),
    .io_ho_input(bc_pe_706_io_ho_input),
    .io_ve_input(bc_pe_706_io_ve_input),
    .io_input_valid(bc_pe_706_io_input_valid),
    .io_iormac(bc_pe_706_io_iormac),
    .io_ve_out(bc_pe_706_io_ve_out),
    .io_ho_out(bc_pe_706_io_ho_out),
    .io_res_out(bc_pe_706_io_res_out)
  );
  bc_pe bc_pe_707 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_707_clock),
    .reset(bc_pe_707_reset),
    .io_ho_input(bc_pe_707_io_ho_input),
    .io_ve_input(bc_pe_707_io_ve_input),
    .io_input_valid(bc_pe_707_io_input_valid),
    .io_iormac(bc_pe_707_io_iormac),
    .io_ve_out(bc_pe_707_io_ve_out),
    .io_ho_out(bc_pe_707_io_ho_out),
    .io_res_out(bc_pe_707_io_res_out)
  );
  bc_pe bc_pe_708 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_708_clock),
    .reset(bc_pe_708_reset),
    .io_ho_input(bc_pe_708_io_ho_input),
    .io_ve_input(bc_pe_708_io_ve_input),
    .io_input_valid(bc_pe_708_io_input_valid),
    .io_iormac(bc_pe_708_io_iormac),
    .io_ve_out(bc_pe_708_io_ve_out),
    .io_ho_out(bc_pe_708_io_ho_out),
    .io_res_out(bc_pe_708_io_res_out)
  );
  bc_pe bc_pe_709 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_709_clock),
    .reset(bc_pe_709_reset),
    .io_ho_input(bc_pe_709_io_ho_input),
    .io_ve_input(bc_pe_709_io_ve_input),
    .io_input_valid(bc_pe_709_io_input_valid),
    .io_iormac(bc_pe_709_io_iormac),
    .io_ve_out(bc_pe_709_io_ve_out),
    .io_ho_out(bc_pe_709_io_ho_out),
    .io_res_out(bc_pe_709_io_res_out)
  );
  bc_pe bc_pe_710 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_710_clock),
    .reset(bc_pe_710_reset),
    .io_ho_input(bc_pe_710_io_ho_input),
    .io_ve_input(bc_pe_710_io_ve_input),
    .io_input_valid(bc_pe_710_io_input_valid),
    .io_iormac(bc_pe_710_io_iormac),
    .io_ve_out(bc_pe_710_io_ve_out),
    .io_ho_out(bc_pe_710_io_ho_out),
    .io_res_out(bc_pe_710_io_res_out)
  );
  bc_pe bc_pe_711 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_711_clock),
    .reset(bc_pe_711_reset),
    .io_ho_input(bc_pe_711_io_ho_input),
    .io_ve_input(bc_pe_711_io_ve_input),
    .io_input_valid(bc_pe_711_io_input_valid),
    .io_iormac(bc_pe_711_io_iormac),
    .io_ve_out(bc_pe_711_io_ve_out),
    .io_ho_out(bc_pe_711_io_ho_out),
    .io_res_out(bc_pe_711_io_res_out)
  );
  bc_pe bc_pe_712 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_712_clock),
    .reset(bc_pe_712_reset),
    .io_ho_input(bc_pe_712_io_ho_input),
    .io_ve_input(bc_pe_712_io_ve_input),
    .io_input_valid(bc_pe_712_io_input_valid),
    .io_iormac(bc_pe_712_io_iormac),
    .io_ve_out(bc_pe_712_io_ve_out),
    .io_ho_out(bc_pe_712_io_ho_out),
    .io_res_out(bc_pe_712_io_res_out)
  );
  bc_pe bc_pe_713 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_713_clock),
    .reset(bc_pe_713_reset),
    .io_ho_input(bc_pe_713_io_ho_input),
    .io_ve_input(bc_pe_713_io_ve_input),
    .io_input_valid(bc_pe_713_io_input_valid),
    .io_iormac(bc_pe_713_io_iormac),
    .io_ve_out(bc_pe_713_io_ve_out),
    .io_ho_out(bc_pe_713_io_ho_out),
    .io_res_out(bc_pe_713_io_res_out)
  );
  bc_pe bc_pe_714 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_714_clock),
    .reset(bc_pe_714_reset),
    .io_ho_input(bc_pe_714_io_ho_input),
    .io_ve_input(bc_pe_714_io_ve_input),
    .io_input_valid(bc_pe_714_io_input_valid),
    .io_iormac(bc_pe_714_io_iormac),
    .io_ve_out(bc_pe_714_io_ve_out),
    .io_ho_out(bc_pe_714_io_ho_out),
    .io_res_out(bc_pe_714_io_res_out)
  );
  bc_pe bc_pe_715 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_715_clock),
    .reset(bc_pe_715_reset),
    .io_ho_input(bc_pe_715_io_ho_input),
    .io_ve_input(bc_pe_715_io_ve_input),
    .io_input_valid(bc_pe_715_io_input_valid),
    .io_iormac(bc_pe_715_io_iormac),
    .io_ve_out(bc_pe_715_io_ve_out),
    .io_ho_out(bc_pe_715_io_ho_out),
    .io_res_out(bc_pe_715_io_res_out)
  );
  bc_pe bc_pe_716 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_716_clock),
    .reset(bc_pe_716_reset),
    .io_ho_input(bc_pe_716_io_ho_input),
    .io_ve_input(bc_pe_716_io_ve_input),
    .io_input_valid(bc_pe_716_io_input_valid),
    .io_iormac(bc_pe_716_io_iormac),
    .io_ve_out(bc_pe_716_io_ve_out),
    .io_ho_out(bc_pe_716_io_ho_out),
    .io_res_out(bc_pe_716_io_res_out)
  );
  bc_pe bc_pe_717 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_717_clock),
    .reset(bc_pe_717_reset),
    .io_ho_input(bc_pe_717_io_ho_input),
    .io_ve_input(bc_pe_717_io_ve_input),
    .io_input_valid(bc_pe_717_io_input_valid),
    .io_iormac(bc_pe_717_io_iormac),
    .io_ve_out(bc_pe_717_io_ve_out),
    .io_ho_out(bc_pe_717_io_ho_out),
    .io_res_out(bc_pe_717_io_res_out)
  );
  bc_pe bc_pe_718 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_718_clock),
    .reset(bc_pe_718_reset),
    .io_ho_input(bc_pe_718_io_ho_input),
    .io_ve_input(bc_pe_718_io_ve_input),
    .io_input_valid(bc_pe_718_io_input_valid),
    .io_iormac(bc_pe_718_io_iormac),
    .io_ve_out(bc_pe_718_io_ve_out),
    .io_ho_out(bc_pe_718_io_ho_out),
    .io_res_out(bc_pe_718_io_res_out)
  );
  bc_pe bc_pe_719 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_719_clock),
    .reset(bc_pe_719_reset),
    .io_ho_input(bc_pe_719_io_ho_input),
    .io_ve_input(bc_pe_719_io_ve_input),
    .io_input_valid(bc_pe_719_io_input_valid),
    .io_iormac(bc_pe_719_io_iormac),
    .io_ve_out(bc_pe_719_io_ve_out),
    .io_ho_out(bc_pe_719_io_ho_out),
    .io_res_out(bc_pe_719_io_res_out)
  );
  bc_pe bc_pe_720 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_720_clock),
    .reset(bc_pe_720_reset),
    .io_ho_input(bc_pe_720_io_ho_input),
    .io_ve_input(bc_pe_720_io_ve_input),
    .io_input_valid(bc_pe_720_io_input_valid),
    .io_iormac(bc_pe_720_io_iormac),
    .io_ve_out(bc_pe_720_io_ve_out),
    .io_ho_out(bc_pe_720_io_ho_out),
    .io_res_out(bc_pe_720_io_res_out)
  );
  bc_pe bc_pe_721 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_721_clock),
    .reset(bc_pe_721_reset),
    .io_ho_input(bc_pe_721_io_ho_input),
    .io_ve_input(bc_pe_721_io_ve_input),
    .io_input_valid(bc_pe_721_io_input_valid),
    .io_iormac(bc_pe_721_io_iormac),
    .io_ve_out(bc_pe_721_io_ve_out),
    .io_ho_out(bc_pe_721_io_ho_out),
    .io_res_out(bc_pe_721_io_res_out)
  );
  bc_pe bc_pe_722 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_722_clock),
    .reset(bc_pe_722_reset),
    .io_ho_input(bc_pe_722_io_ho_input),
    .io_ve_input(bc_pe_722_io_ve_input),
    .io_input_valid(bc_pe_722_io_input_valid),
    .io_iormac(bc_pe_722_io_iormac),
    .io_ve_out(bc_pe_722_io_ve_out),
    .io_ho_out(bc_pe_722_io_ho_out),
    .io_res_out(bc_pe_722_io_res_out)
  );
  bc_pe bc_pe_723 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_723_clock),
    .reset(bc_pe_723_reset),
    .io_ho_input(bc_pe_723_io_ho_input),
    .io_ve_input(bc_pe_723_io_ve_input),
    .io_input_valid(bc_pe_723_io_input_valid),
    .io_iormac(bc_pe_723_io_iormac),
    .io_ve_out(bc_pe_723_io_ve_out),
    .io_ho_out(bc_pe_723_io_ho_out),
    .io_res_out(bc_pe_723_io_res_out)
  );
  bc_pe bc_pe_724 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_724_clock),
    .reset(bc_pe_724_reset),
    .io_ho_input(bc_pe_724_io_ho_input),
    .io_ve_input(bc_pe_724_io_ve_input),
    .io_input_valid(bc_pe_724_io_input_valid),
    .io_iormac(bc_pe_724_io_iormac),
    .io_ve_out(bc_pe_724_io_ve_out),
    .io_ho_out(bc_pe_724_io_ho_out),
    .io_res_out(bc_pe_724_io_res_out)
  );
  bc_pe bc_pe_725 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_725_clock),
    .reset(bc_pe_725_reset),
    .io_ho_input(bc_pe_725_io_ho_input),
    .io_ve_input(bc_pe_725_io_ve_input),
    .io_input_valid(bc_pe_725_io_input_valid),
    .io_iormac(bc_pe_725_io_iormac),
    .io_ve_out(bc_pe_725_io_ve_out),
    .io_ho_out(bc_pe_725_io_ho_out),
    .io_res_out(bc_pe_725_io_res_out)
  );
  bc_pe bc_pe_726 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_726_clock),
    .reset(bc_pe_726_reset),
    .io_ho_input(bc_pe_726_io_ho_input),
    .io_ve_input(bc_pe_726_io_ve_input),
    .io_input_valid(bc_pe_726_io_input_valid),
    .io_iormac(bc_pe_726_io_iormac),
    .io_ve_out(bc_pe_726_io_ve_out),
    .io_ho_out(bc_pe_726_io_ho_out),
    .io_res_out(bc_pe_726_io_res_out)
  );
  bc_pe bc_pe_727 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_727_clock),
    .reset(bc_pe_727_reset),
    .io_ho_input(bc_pe_727_io_ho_input),
    .io_ve_input(bc_pe_727_io_ve_input),
    .io_input_valid(bc_pe_727_io_input_valid),
    .io_iormac(bc_pe_727_io_iormac),
    .io_ve_out(bc_pe_727_io_ve_out),
    .io_ho_out(bc_pe_727_io_ho_out),
    .io_res_out(bc_pe_727_io_res_out)
  );
  bc_pe bc_pe_728 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_728_clock),
    .reset(bc_pe_728_reset),
    .io_ho_input(bc_pe_728_io_ho_input),
    .io_ve_input(bc_pe_728_io_ve_input),
    .io_input_valid(bc_pe_728_io_input_valid),
    .io_iormac(bc_pe_728_io_iormac),
    .io_ve_out(bc_pe_728_io_ve_out),
    .io_ho_out(bc_pe_728_io_ho_out),
    .io_res_out(bc_pe_728_io_res_out)
  );
  bc_pe bc_pe_729 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_729_clock),
    .reset(bc_pe_729_reset),
    .io_ho_input(bc_pe_729_io_ho_input),
    .io_ve_input(bc_pe_729_io_ve_input),
    .io_input_valid(bc_pe_729_io_input_valid),
    .io_iormac(bc_pe_729_io_iormac),
    .io_ve_out(bc_pe_729_io_ve_out),
    .io_ho_out(bc_pe_729_io_ho_out),
    .io_res_out(bc_pe_729_io_res_out)
  );
  bc_pe bc_pe_730 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_730_clock),
    .reset(bc_pe_730_reset),
    .io_ho_input(bc_pe_730_io_ho_input),
    .io_ve_input(bc_pe_730_io_ve_input),
    .io_input_valid(bc_pe_730_io_input_valid),
    .io_iormac(bc_pe_730_io_iormac),
    .io_ve_out(bc_pe_730_io_ve_out),
    .io_ho_out(bc_pe_730_io_ho_out),
    .io_res_out(bc_pe_730_io_res_out)
  );
  bc_pe bc_pe_731 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_731_clock),
    .reset(bc_pe_731_reset),
    .io_ho_input(bc_pe_731_io_ho_input),
    .io_ve_input(bc_pe_731_io_ve_input),
    .io_input_valid(bc_pe_731_io_input_valid),
    .io_iormac(bc_pe_731_io_iormac),
    .io_ve_out(bc_pe_731_io_ve_out),
    .io_ho_out(bc_pe_731_io_ho_out),
    .io_res_out(bc_pe_731_io_res_out)
  );
  bc_pe bc_pe_732 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_732_clock),
    .reset(bc_pe_732_reset),
    .io_ho_input(bc_pe_732_io_ho_input),
    .io_ve_input(bc_pe_732_io_ve_input),
    .io_input_valid(bc_pe_732_io_input_valid),
    .io_iormac(bc_pe_732_io_iormac),
    .io_ve_out(bc_pe_732_io_ve_out),
    .io_ho_out(bc_pe_732_io_ho_out),
    .io_res_out(bc_pe_732_io_res_out)
  );
  bc_pe bc_pe_733 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_733_clock),
    .reset(bc_pe_733_reset),
    .io_ho_input(bc_pe_733_io_ho_input),
    .io_ve_input(bc_pe_733_io_ve_input),
    .io_input_valid(bc_pe_733_io_input_valid),
    .io_iormac(bc_pe_733_io_iormac),
    .io_ve_out(bc_pe_733_io_ve_out),
    .io_ho_out(bc_pe_733_io_ho_out),
    .io_res_out(bc_pe_733_io_res_out)
  );
  bc_pe bc_pe_734 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_734_clock),
    .reset(bc_pe_734_reset),
    .io_ho_input(bc_pe_734_io_ho_input),
    .io_ve_input(bc_pe_734_io_ve_input),
    .io_input_valid(bc_pe_734_io_input_valid),
    .io_iormac(bc_pe_734_io_iormac),
    .io_ve_out(bc_pe_734_io_ve_out),
    .io_ho_out(bc_pe_734_io_ho_out),
    .io_res_out(bc_pe_734_io_res_out)
  );
  bc_pe bc_pe_735 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_735_clock),
    .reset(bc_pe_735_reset),
    .io_ho_input(bc_pe_735_io_ho_input),
    .io_ve_input(bc_pe_735_io_ve_input),
    .io_input_valid(bc_pe_735_io_input_valid),
    .io_iormac(bc_pe_735_io_iormac),
    .io_ve_out(bc_pe_735_io_ve_out),
    .io_ho_out(bc_pe_735_io_ho_out),
    .io_res_out(bc_pe_735_io_res_out)
  );
  bc_pe bc_pe_736 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_736_clock),
    .reset(bc_pe_736_reset),
    .io_ho_input(bc_pe_736_io_ho_input),
    .io_ve_input(bc_pe_736_io_ve_input),
    .io_input_valid(bc_pe_736_io_input_valid),
    .io_iormac(bc_pe_736_io_iormac),
    .io_ve_out(bc_pe_736_io_ve_out),
    .io_ho_out(bc_pe_736_io_ho_out),
    .io_res_out(bc_pe_736_io_res_out)
  );
  bc_pe bc_pe_737 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_737_clock),
    .reset(bc_pe_737_reset),
    .io_ho_input(bc_pe_737_io_ho_input),
    .io_ve_input(bc_pe_737_io_ve_input),
    .io_input_valid(bc_pe_737_io_input_valid),
    .io_iormac(bc_pe_737_io_iormac),
    .io_ve_out(bc_pe_737_io_ve_out),
    .io_ho_out(bc_pe_737_io_ho_out),
    .io_res_out(bc_pe_737_io_res_out)
  );
  bc_pe bc_pe_738 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_738_clock),
    .reset(bc_pe_738_reset),
    .io_ho_input(bc_pe_738_io_ho_input),
    .io_ve_input(bc_pe_738_io_ve_input),
    .io_input_valid(bc_pe_738_io_input_valid),
    .io_iormac(bc_pe_738_io_iormac),
    .io_ve_out(bc_pe_738_io_ve_out),
    .io_ho_out(bc_pe_738_io_ho_out),
    .io_res_out(bc_pe_738_io_res_out)
  );
  bc_pe bc_pe_739 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_739_clock),
    .reset(bc_pe_739_reset),
    .io_ho_input(bc_pe_739_io_ho_input),
    .io_ve_input(bc_pe_739_io_ve_input),
    .io_input_valid(bc_pe_739_io_input_valid),
    .io_iormac(bc_pe_739_io_iormac),
    .io_ve_out(bc_pe_739_io_ve_out),
    .io_ho_out(bc_pe_739_io_ho_out),
    .io_res_out(bc_pe_739_io_res_out)
  );
  bc_pe bc_pe_740 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_740_clock),
    .reset(bc_pe_740_reset),
    .io_ho_input(bc_pe_740_io_ho_input),
    .io_ve_input(bc_pe_740_io_ve_input),
    .io_input_valid(bc_pe_740_io_input_valid),
    .io_iormac(bc_pe_740_io_iormac),
    .io_ve_out(bc_pe_740_io_ve_out),
    .io_ho_out(bc_pe_740_io_ho_out),
    .io_res_out(bc_pe_740_io_res_out)
  );
  bc_pe bc_pe_741 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_741_clock),
    .reset(bc_pe_741_reset),
    .io_ho_input(bc_pe_741_io_ho_input),
    .io_ve_input(bc_pe_741_io_ve_input),
    .io_input_valid(bc_pe_741_io_input_valid),
    .io_iormac(bc_pe_741_io_iormac),
    .io_ve_out(bc_pe_741_io_ve_out),
    .io_ho_out(bc_pe_741_io_ho_out),
    .io_res_out(bc_pe_741_io_res_out)
  );
  bc_pe bc_pe_742 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_742_clock),
    .reset(bc_pe_742_reset),
    .io_ho_input(bc_pe_742_io_ho_input),
    .io_ve_input(bc_pe_742_io_ve_input),
    .io_input_valid(bc_pe_742_io_input_valid),
    .io_iormac(bc_pe_742_io_iormac),
    .io_ve_out(bc_pe_742_io_ve_out),
    .io_ho_out(bc_pe_742_io_ho_out),
    .io_res_out(bc_pe_742_io_res_out)
  );
  bc_pe bc_pe_743 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_743_clock),
    .reset(bc_pe_743_reset),
    .io_ho_input(bc_pe_743_io_ho_input),
    .io_ve_input(bc_pe_743_io_ve_input),
    .io_input_valid(bc_pe_743_io_input_valid),
    .io_iormac(bc_pe_743_io_iormac),
    .io_ve_out(bc_pe_743_io_ve_out),
    .io_ho_out(bc_pe_743_io_ho_out),
    .io_res_out(bc_pe_743_io_res_out)
  );
  bc_pe bc_pe_744 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_744_clock),
    .reset(bc_pe_744_reset),
    .io_ho_input(bc_pe_744_io_ho_input),
    .io_ve_input(bc_pe_744_io_ve_input),
    .io_input_valid(bc_pe_744_io_input_valid),
    .io_iormac(bc_pe_744_io_iormac),
    .io_ve_out(bc_pe_744_io_ve_out),
    .io_ho_out(bc_pe_744_io_ho_out),
    .io_res_out(bc_pe_744_io_res_out)
  );
  bc_pe bc_pe_745 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_745_clock),
    .reset(bc_pe_745_reset),
    .io_ho_input(bc_pe_745_io_ho_input),
    .io_ve_input(bc_pe_745_io_ve_input),
    .io_input_valid(bc_pe_745_io_input_valid),
    .io_iormac(bc_pe_745_io_iormac),
    .io_ve_out(bc_pe_745_io_ve_out),
    .io_ho_out(bc_pe_745_io_ho_out),
    .io_res_out(bc_pe_745_io_res_out)
  );
  bc_pe bc_pe_746 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_746_clock),
    .reset(bc_pe_746_reset),
    .io_ho_input(bc_pe_746_io_ho_input),
    .io_ve_input(bc_pe_746_io_ve_input),
    .io_input_valid(bc_pe_746_io_input_valid),
    .io_iormac(bc_pe_746_io_iormac),
    .io_ve_out(bc_pe_746_io_ve_out),
    .io_ho_out(bc_pe_746_io_ho_out),
    .io_res_out(bc_pe_746_io_res_out)
  );
  bc_pe bc_pe_747 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_747_clock),
    .reset(bc_pe_747_reset),
    .io_ho_input(bc_pe_747_io_ho_input),
    .io_ve_input(bc_pe_747_io_ve_input),
    .io_input_valid(bc_pe_747_io_input_valid),
    .io_iormac(bc_pe_747_io_iormac),
    .io_ve_out(bc_pe_747_io_ve_out),
    .io_ho_out(bc_pe_747_io_ho_out),
    .io_res_out(bc_pe_747_io_res_out)
  );
  bc_pe bc_pe_748 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_748_clock),
    .reset(bc_pe_748_reset),
    .io_ho_input(bc_pe_748_io_ho_input),
    .io_ve_input(bc_pe_748_io_ve_input),
    .io_input_valid(bc_pe_748_io_input_valid),
    .io_iormac(bc_pe_748_io_iormac),
    .io_ve_out(bc_pe_748_io_ve_out),
    .io_ho_out(bc_pe_748_io_ho_out),
    .io_res_out(bc_pe_748_io_res_out)
  );
  bc_pe bc_pe_749 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_749_clock),
    .reset(bc_pe_749_reset),
    .io_ho_input(bc_pe_749_io_ho_input),
    .io_ve_input(bc_pe_749_io_ve_input),
    .io_input_valid(bc_pe_749_io_input_valid),
    .io_iormac(bc_pe_749_io_iormac),
    .io_ve_out(bc_pe_749_io_ve_out),
    .io_ho_out(bc_pe_749_io_ho_out),
    .io_res_out(bc_pe_749_io_res_out)
  );
  bc_pe bc_pe_750 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_750_clock),
    .reset(bc_pe_750_reset),
    .io_ho_input(bc_pe_750_io_ho_input),
    .io_ve_input(bc_pe_750_io_ve_input),
    .io_input_valid(bc_pe_750_io_input_valid),
    .io_iormac(bc_pe_750_io_iormac),
    .io_ve_out(bc_pe_750_io_ve_out),
    .io_ho_out(bc_pe_750_io_ho_out),
    .io_res_out(bc_pe_750_io_res_out)
  );
  bc_pe bc_pe_751 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_751_clock),
    .reset(bc_pe_751_reset),
    .io_ho_input(bc_pe_751_io_ho_input),
    .io_ve_input(bc_pe_751_io_ve_input),
    .io_input_valid(bc_pe_751_io_input_valid),
    .io_iormac(bc_pe_751_io_iormac),
    .io_ve_out(bc_pe_751_io_ve_out),
    .io_ho_out(bc_pe_751_io_ho_out),
    .io_res_out(bc_pe_751_io_res_out)
  );
  bc_pe bc_pe_752 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_752_clock),
    .reset(bc_pe_752_reset),
    .io_ho_input(bc_pe_752_io_ho_input),
    .io_ve_input(bc_pe_752_io_ve_input),
    .io_input_valid(bc_pe_752_io_input_valid),
    .io_iormac(bc_pe_752_io_iormac),
    .io_ve_out(bc_pe_752_io_ve_out),
    .io_ho_out(bc_pe_752_io_ho_out),
    .io_res_out(bc_pe_752_io_res_out)
  );
  bc_pe bc_pe_753 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_753_clock),
    .reset(bc_pe_753_reset),
    .io_ho_input(bc_pe_753_io_ho_input),
    .io_ve_input(bc_pe_753_io_ve_input),
    .io_input_valid(bc_pe_753_io_input_valid),
    .io_iormac(bc_pe_753_io_iormac),
    .io_ve_out(bc_pe_753_io_ve_out),
    .io_ho_out(bc_pe_753_io_ho_out),
    .io_res_out(bc_pe_753_io_res_out)
  );
  bc_pe bc_pe_754 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_754_clock),
    .reset(bc_pe_754_reset),
    .io_ho_input(bc_pe_754_io_ho_input),
    .io_ve_input(bc_pe_754_io_ve_input),
    .io_input_valid(bc_pe_754_io_input_valid),
    .io_iormac(bc_pe_754_io_iormac),
    .io_ve_out(bc_pe_754_io_ve_out),
    .io_ho_out(bc_pe_754_io_ho_out),
    .io_res_out(bc_pe_754_io_res_out)
  );
  bc_pe bc_pe_755 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_755_clock),
    .reset(bc_pe_755_reset),
    .io_ho_input(bc_pe_755_io_ho_input),
    .io_ve_input(bc_pe_755_io_ve_input),
    .io_input_valid(bc_pe_755_io_input_valid),
    .io_iormac(bc_pe_755_io_iormac),
    .io_ve_out(bc_pe_755_io_ve_out),
    .io_ho_out(bc_pe_755_io_ho_out),
    .io_res_out(bc_pe_755_io_res_out)
  );
  bc_pe bc_pe_756 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_756_clock),
    .reset(bc_pe_756_reset),
    .io_ho_input(bc_pe_756_io_ho_input),
    .io_ve_input(bc_pe_756_io_ve_input),
    .io_input_valid(bc_pe_756_io_input_valid),
    .io_iormac(bc_pe_756_io_iormac),
    .io_ve_out(bc_pe_756_io_ve_out),
    .io_ho_out(bc_pe_756_io_ho_out),
    .io_res_out(bc_pe_756_io_res_out)
  );
  bc_pe bc_pe_757 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_757_clock),
    .reset(bc_pe_757_reset),
    .io_ho_input(bc_pe_757_io_ho_input),
    .io_ve_input(bc_pe_757_io_ve_input),
    .io_input_valid(bc_pe_757_io_input_valid),
    .io_iormac(bc_pe_757_io_iormac),
    .io_ve_out(bc_pe_757_io_ve_out),
    .io_ho_out(bc_pe_757_io_ho_out),
    .io_res_out(bc_pe_757_io_res_out)
  );
  bc_pe bc_pe_758 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_758_clock),
    .reset(bc_pe_758_reset),
    .io_ho_input(bc_pe_758_io_ho_input),
    .io_ve_input(bc_pe_758_io_ve_input),
    .io_input_valid(bc_pe_758_io_input_valid),
    .io_iormac(bc_pe_758_io_iormac),
    .io_ve_out(bc_pe_758_io_ve_out),
    .io_ho_out(bc_pe_758_io_ho_out),
    .io_res_out(bc_pe_758_io_res_out)
  );
  bc_pe bc_pe_759 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_759_clock),
    .reset(bc_pe_759_reset),
    .io_ho_input(bc_pe_759_io_ho_input),
    .io_ve_input(bc_pe_759_io_ve_input),
    .io_input_valid(bc_pe_759_io_input_valid),
    .io_iormac(bc_pe_759_io_iormac),
    .io_ve_out(bc_pe_759_io_ve_out),
    .io_ho_out(bc_pe_759_io_ho_out),
    .io_res_out(bc_pe_759_io_res_out)
  );
  bc_pe bc_pe_760 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_760_clock),
    .reset(bc_pe_760_reset),
    .io_ho_input(bc_pe_760_io_ho_input),
    .io_ve_input(bc_pe_760_io_ve_input),
    .io_input_valid(bc_pe_760_io_input_valid),
    .io_iormac(bc_pe_760_io_iormac),
    .io_ve_out(bc_pe_760_io_ve_out),
    .io_ho_out(bc_pe_760_io_ho_out),
    .io_res_out(bc_pe_760_io_res_out)
  );
  bc_pe bc_pe_761 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_761_clock),
    .reset(bc_pe_761_reset),
    .io_ho_input(bc_pe_761_io_ho_input),
    .io_ve_input(bc_pe_761_io_ve_input),
    .io_input_valid(bc_pe_761_io_input_valid),
    .io_iormac(bc_pe_761_io_iormac),
    .io_ve_out(bc_pe_761_io_ve_out),
    .io_ho_out(bc_pe_761_io_ho_out),
    .io_res_out(bc_pe_761_io_res_out)
  );
  bc_pe bc_pe_762 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_762_clock),
    .reset(bc_pe_762_reset),
    .io_ho_input(bc_pe_762_io_ho_input),
    .io_ve_input(bc_pe_762_io_ve_input),
    .io_input_valid(bc_pe_762_io_input_valid),
    .io_iormac(bc_pe_762_io_iormac),
    .io_ve_out(bc_pe_762_io_ve_out),
    .io_ho_out(bc_pe_762_io_ho_out),
    .io_res_out(bc_pe_762_io_res_out)
  );
  bc_pe bc_pe_763 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_763_clock),
    .reset(bc_pe_763_reset),
    .io_ho_input(bc_pe_763_io_ho_input),
    .io_ve_input(bc_pe_763_io_ve_input),
    .io_input_valid(bc_pe_763_io_input_valid),
    .io_iormac(bc_pe_763_io_iormac),
    .io_ve_out(bc_pe_763_io_ve_out),
    .io_ho_out(bc_pe_763_io_ho_out),
    .io_res_out(bc_pe_763_io_res_out)
  );
  bc_pe bc_pe_764 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_764_clock),
    .reset(bc_pe_764_reset),
    .io_ho_input(bc_pe_764_io_ho_input),
    .io_ve_input(bc_pe_764_io_ve_input),
    .io_input_valid(bc_pe_764_io_input_valid),
    .io_iormac(bc_pe_764_io_iormac),
    .io_ve_out(bc_pe_764_io_ve_out),
    .io_ho_out(bc_pe_764_io_ho_out),
    .io_res_out(bc_pe_764_io_res_out)
  );
  bc_pe bc_pe_765 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_765_clock),
    .reset(bc_pe_765_reset),
    .io_ho_input(bc_pe_765_io_ho_input),
    .io_ve_input(bc_pe_765_io_ve_input),
    .io_input_valid(bc_pe_765_io_input_valid),
    .io_iormac(bc_pe_765_io_iormac),
    .io_ve_out(bc_pe_765_io_ve_out),
    .io_ho_out(bc_pe_765_io_ho_out),
    .io_res_out(bc_pe_765_io_res_out)
  );
  bc_pe bc_pe_766 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_766_clock),
    .reset(bc_pe_766_reset),
    .io_ho_input(bc_pe_766_io_ho_input),
    .io_ve_input(bc_pe_766_io_ve_input),
    .io_input_valid(bc_pe_766_io_input_valid),
    .io_iormac(bc_pe_766_io_iormac),
    .io_ve_out(bc_pe_766_io_ve_out),
    .io_ho_out(bc_pe_766_io_ho_out),
    .io_res_out(bc_pe_766_io_res_out)
  );
  bc_pe bc_pe_767 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_767_clock),
    .reset(bc_pe_767_reset),
    .io_ho_input(bc_pe_767_io_ho_input),
    .io_ve_input(bc_pe_767_io_ve_input),
    .io_input_valid(bc_pe_767_io_input_valid),
    .io_iormac(bc_pe_767_io_iormac),
    .io_ve_out(bc_pe_767_io_ve_out),
    .io_ho_out(bc_pe_767_io_ho_out),
    .io_res_out(bc_pe_767_io_res_out)
  );
  bc_pe bc_pe_768 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_768_clock),
    .reset(bc_pe_768_reset),
    .io_ho_input(bc_pe_768_io_ho_input),
    .io_ve_input(bc_pe_768_io_ve_input),
    .io_input_valid(bc_pe_768_io_input_valid),
    .io_iormac(bc_pe_768_io_iormac),
    .io_ve_out(bc_pe_768_io_ve_out),
    .io_ho_out(bc_pe_768_io_ho_out),
    .io_res_out(bc_pe_768_io_res_out)
  );
  bc_pe bc_pe_769 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_769_clock),
    .reset(bc_pe_769_reset),
    .io_ho_input(bc_pe_769_io_ho_input),
    .io_ve_input(bc_pe_769_io_ve_input),
    .io_input_valid(bc_pe_769_io_input_valid),
    .io_iormac(bc_pe_769_io_iormac),
    .io_ve_out(bc_pe_769_io_ve_out),
    .io_ho_out(bc_pe_769_io_ho_out),
    .io_res_out(bc_pe_769_io_res_out)
  );
  bc_pe bc_pe_770 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_770_clock),
    .reset(bc_pe_770_reset),
    .io_ho_input(bc_pe_770_io_ho_input),
    .io_ve_input(bc_pe_770_io_ve_input),
    .io_input_valid(bc_pe_770_io_input_valid),
    .io_iormac(bc_pe_770_io_iormac),
    .io_ve_out(bc_pe_770_io_ve_out),
    .io_ho_out(bc_pe_770_io_ho_out),
    .io_res_out(bc_pe_770_io_res_out)
  );
  bc_pe bc_pe_771 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_771_clock),
    .reset(bc_pe_771_reset),
    .io_ho_input(bc_pe_771_io_ho_input),
    .io_ve_input(bc_pe_771_io_ve_input),
    .io_input_valid(bc_pe_771_io_input_valid),
    .io_iormac(bc_pe_771_io_iormac),
    .io_ve_out(bc_pe_771_io_ve_out),
    .io_ho_out(bc_pe_771_io_ho_out),
    .io_res_out(bc_pe_771_io_res_out)
  );
  bc_pe bc_pe_772 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_772_clock),
    .reset(bc_pe_772_reset),
    .io_ho_input(bc_pe_772_io_ho_input),
    .io_ve_input(bc_pe_772_io_ve_input),
    .io_input_valid(bc_pe_772_io_input_valid),
    .io_iormac(bc_pe_772_io_iormac),
    .io_ve_out(bc_pe_772_io_ve_out),
    .io_ho_out(bc_pe_772_io_ho_out),
    .io_res_out(bc_pe_772_io_res_out)
  );
  bc_pe bc_pe_773 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_773_clock),
    .reset(bc_pe_773_reset),
    .io_ho_input(bc_pe_773_io_ho_input),
    .io_ve_input(bc_pe_773_io_ve_input),
    .io_input_valid(bc_pe_773_io_input_valid),
    .io_iormac(bc_pe_773_io_iormac),
    .io_ve_out(bc_pe_773_io_ve_out),
    .io_ho_out(bc_pe_773_io_ho_out),
    .io_res_out(bc_pe_773_io_res_out)
  );
  bc_pe bc_pe_774 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_774_clock),
    .reset(bc_pe_774_reset),
    .io_ho_input(bc_pe_774_io_ho_input),
    .io_ve_input(bc_pe_774_io_ve_input),
    .io_input_valid(bc_pe_774_io_input_valid),
    .io_iormac(bc_pe_774_io_iormac),
    .io_ve_out(bc_pe_774_io_ve_out),
    .io_ho_out(bc_pe_774_io_ho_out),
    .io_res_out(bc_pe_774_io_res_out)
  );
  bc_pe bc_pe_775 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_775_clock),
    .reset(bc_pe_775_reset),
    .io_ho_input(bc_pe_775_io_ho_input),
    .io_ve_input(bc_pe_775_io_ve_input),
    .io_input_valid(bc_pe_775_io_input_valid),
    .io_iormac(bc_pe_775_io_iormac),
    .io_ve_out(bc_pe_775_io_ve_out),
    .io_ho_out(bc_pe_775_io_ho_out),
    .io_res_out(bc_pe_775_io_res_out)
  );
  bc_pe bc_pe_776 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_776_clock),
    .reset(bc_pe_776_reset),
    .io_ho_input(bc_pe_776_io_ho_input),
    .io_ve_input(bc_pe_776_io_ve_input),
    .io_input_valid(bc_pe_776_io_input_valid),
    .io_iormac(bc_pe_776_io_iormac),
    .io_ve_out(bc_pe_776_io_ve_out),
    .io_ho_out(bc_pe_776_io_ho_out),
    .io_res_out(bc_pe_776_io_res_out)
  );
  bc_pe bc_pe_777 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_777_clock),
    .reset(bc_pe_777_reset),
    .io_ho_input(bc_pe_777_io_ho_input),
    .io_ve_input(bc_pe_777_io_ve_input),
    .io_input_valid(bc_pe_777_io_input_valid),
    .io_iormac(bc_pe_777_io_iormac),
    .io_ve_out(bc_pe_777_io_ve_out),
    .io_ho_out(bc_pe_777_io_ho_out),
    .io_res_out(bc_pe_777_io_res_out)
  );
  bc_pe bc_pe_778 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_778_clock),
    .reset(bc_pe_778_reset),
    .io_ho_input(bc_pe_778_io_ho_input),
    .io_ve_input(bc_pe_778_io_ve_input),
    .io_input_valid(bc_pe_778_io_input_valid),
    .io_iormac(bc_pe_778_io_iormac),
    .io_ve_out(bc_pe_778_io_ve_out),
    .io_ho_out(bc_pe_778_io_ho_out),
    .io_res_out(bc_pe_778_io_res_out)
  );
  bc_pe bc_pe_779 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_779_clock),
    .reset(bc_pe_779_reset),
    .io_ho_input(bc_pe_779_io_ho_input),
    .io_ve_input(bc_pe_779_io_ve_input),
    .io_input_valid(bc_pe_779_io_input_valid),
    .io_iormac(bc_pe_779_io_iormac),
    .io_ve_out(bc_pe_779_io_ve_out),
    .io_ho_out(bc_pe_779_io_ho_out),
    .io_res_out(bc_pe_779_io_res_out)
  );
  bc_pe bc_pe_780 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_780_clock),
    .reset(bc_pe_780_reset),
    .io_ho_input(bc_pe_780_io_ho_input),
    .io_ve_input(bc_pe_780_io_ve_input),
    .io_input_valid(bc_pe_780_io_input_valid),
    .io_iormac(bc_pe_780_io_iormac),
    .io_ve_out(bc_pe_780_io_ve_out),
    .io_ho_out(bc_pe_780_io_ho_out),
    .io_res_out(bc_pe_780_io_res_out)
  );
  bc_pe bc_pe_781 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_781_clock),
    .reset(bc_pe_781_reset),
    .io_ho_input(bc_pe_781_io_ho_input),
    .io_ve_input(bc_pe_781_io_ve_input),
    .io_input_valid(bc_pe_781_io_input_valid),
    .io_iormac(bc_pe_781_io_iormac),
    .io_ve_out(bc_pe_781_io_ve_out),
    .io_ho_out(bc_pe_781_io_ho_out),
    .io_res_out(bc_pe_781_io_res_out)
  );
  bc_pe bc_pe_782 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_782_clock),
    .reset(bc_pe_782_reset),
    .io_ho_input(bc_pe_782_io_ho_input),
    .io_ve_input(bc_pe_782_io_ve_input),
    .io_input_valid(bc_pe_782_io_input_valid),
    .io_iormac(bc_pe_782_io_iormac),
    .io_ve_out(bc_pe_782_io_ve_out),
    .io_ho_out(bc_pe_782_io_ho_out),
    .io_res_out(bc_pe_782_io_res_out)
  );
  bc_pe bc_pe_783 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_783_clock),
    .reset(bc_pe_783_reset),
    .io_ho_input(bc_pe_783_io_ho_input),
    .io_ve_input(bc_pe_783_io_ve_input),
    .io_input_valid(bc_pe_783_io_input_valid),
    .io_iormac(bc_pe_783_io_iormac),
    .io_ve_out(bc_pe_783_io_ve_out),
    .io_ho_out(bc_pe_783_io_ho_out),
    .io_res_out(bc_pe_783_io_res_out)
  );
  bc_pe bc_pe_784 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_784_clock),
    .reset(bc_pe_784_reset),
    .io_ho_input(bc_pe_784_io_ho_input),
    .io_ve_input(bc_pe_784_io_ve_input),
    .io_input_valid(bc_pe_784_io_input_valid),
    .io_iormac(bc_pe_784_io_iormac),
    .io_ve_out(bc_pe_784_io_ve_out),
    .io_ho_out(bc_pe_784_io_ho_out),
    .io_res_out(bc_pe_784_io_res_out)
  );
  bc_pe bc_pe_785 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_785_clock),
    .reset(bc_pe_785_reset),
    .io_ho_input(bc_pe_785_io_ho_input),
    .io_ve_input(bc_pe_785_io_ve_input),
    .io_input_valid(bc_pe_785_io_input_valid),
    .io_iormac(bc_pe_785_io_iormac),
    .io_ve_out(bc_pe_785_io_ve_out),
    .io_ho_out(bc_pe_785_io_ho_out),
    .io_res_out(bc_pe_785_io_res_out)
  );
  bc_pe bc_pe_786 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_786_clock),
    .reset(bc_pe_786_reset),
    .io_ho_input(bc_pe_786_io_ho_input),
    .io_ve_input(bc_pe_786_io_ve_input),
    .io_input_valid(bc_pe_786_io_input_valid),
    .io_iormac(bc_pe_786_io_iormac),
    .io_ve_out(bc_pe_786_io_ve_out),
    .io_ho_out(bc_pe_786_io_ho_out),
    .io_res_out(bc_pe_786_io_res_out)
  );
  bc_pe bc_pe_787 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_787_clock),
    .reset(bc_pe_787_reset),
    .io_ho_input(bc_pe_787_io_ho_input),
    .io_ve_input(bc_pe_787_io_ve_input),
    .io_input_valid(bc_pe_787_io_input_valid),
    .io_iormac(bc_pe_787_io_iormac),
    .io_ve_out(bc_pe_787_io_ve_out),
    .io_ho_out(bc_pe_787_io_ho_out),
    .io_res_out(bc_pe_787_io_res_out)
  );
  bc_pe bc_pe_788 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_788_clock),
    .reset(bc_pe_788_reset),
    .io_ho_input(bc_pe_788_io_ho_input),
    .io_ve_input(bc_pe_788_io_ve_input),
    .io_input_valid(bc_pe_788_io_input_valid),
    .io_iormac(bc_pe_788_io_iormac),
    .io_ve_out(bc_pe_788_io_ve_out),
    .io_ho_out(bc_pe_788_io_ho_out),
    .io_res_out(bc_pe_788_io_res_out)
  );
  bc_pe bc_pe_789 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_789_clock),
    .reset(bc_pe_789_reset),
    .io_ho_input(bc_pe_789_io_ho_input),
    .io_ve_input(bc_pe_789_io_ve_input),
    .io_input_valid(bc_pe_789_io_input_valid),
    .io_iormac(bc_pe_789_io_iormac),
    .io_ve_out(bc_pe_789_io_ve_out),
    .io_ho_out(bc_pe_789_io_ho_out),
    .io_res_out(bc_pe_789_io_res_out)
  );
  bc_pe bc_pe_790 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_790_clock),
    .reset(bc_pe_790_reset),
    .io_ho_input(bc_pe_790_io_ho_input),
    .io_ve_input(bc_pe_790_io_ve_input),
    .io_input_valid(bc_pe_790_io_input_valid),
    .io_iormac(bc_pe_790_io_iormac),
    .io_ve_out(bc_pe_790_io_ve_out),
    .io_ho_out(bc_pe_790_io_ho_out),
    .io_res_out(bc_pe_790_io_res_out)
  );
  bc_pe bc_pe_791 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_791_clock),
    .reset(bc_pe_791_reset),
    .io_ho_input(bc_pe_791_io_ho_input),
    .io_ve_input(bc_pe_791_io_ve_input),
    .io_input_valid(bc_pe_791_io_input_valid),
    .io_iormac(bc_pe_791_io_iormac),
    .io_ve_out(bc_pe_791_io_ve_out),
    .io_ho_out(bc_pe_791_io_ho_out),
    .io_res_out(bc_pe_791_io_res_out)
  );
  bc_pe bc_pe_792 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_792_clock),
    .reset(bc_pe_792_reset),
    .io_ho_input(bc_pe_792_io_ho_input),
    .io_ve_input(bc_pe_792_io_ve_input),
    .io_input_valid(bc_pe_792_io_input_valid),
    .io_iormac(bc_pe_792_io_iormac),
    .io_ve_out(bc_pe_792_io_ve_out),
    .io_ho_out(bc_pe_792_io_ho_out),
    .io_res_out(bc_pe_792_io_res_out)
  );
  bc_pe bc_pe_793 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_793_clock),
    .reset(bc_pe_793_reset),
    .io_ho_input(bc_pe_793_io_ho_input),
    .io_ve_input(bc_pe_793_io_ve_input),
    .io_input_valid(bc_pe_793_io_input_valid),
    .io_iormac(bc_pe_793_io_iormac),
    .io_ve_out(bc_pe_793_io_ve_out),
    .io_ho_out(bc_pe_793_io_ho_out),
    .io_res_out(bc_pe_793_io_res_out)
  );
  bc_pe bc_pe_794 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_794_clock),
    .reset(bc_pe_794_reset),
    .io_ho_input(bc_pe_794_io_ho_input),
    .io_ve_input(bc_pe_794_io_ve_input),
    .io_input_valid(bc_pe_794_io_input_valid),
    .io_iormac(bc_pe_794_io_iormac),
    .io_ve_out(bc_pe_794_io_ve_out),
    .io_ho_out(bc_pe_794_io_ho_out),
    .io_res_out(bc_pe_794_io_res_out)
  );
  bc_pe bc_pe_795 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_795_clock),
    .reset(bc_pe_795_reset),
    .io_ho_input(bc_pe_795_io_ho_input),
    .io_ve_input(bc_pe_795_io_ve_input),
    .io_input_valid(bc_pe_795_io_input_valid),
    .io_iormac(bc_pe_795_io_iormac),
    .io_ve_out(bc_pe_795_io_ve_out),
    .io_ho_out(bc_pe_795_io_ho_out),
    .io_res_out(bc_pe_795_io_res_out)
  );
  bc_pe bc_pe_796 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_796_clock),
    .reset(bc_pe_796_reset),
    .io_ho_input(bc_pe_796_io_ho_input),
    .io_ve_input(bc_pe_796_io_ve_input),
    .io_input_valid(bc_pe_796_io_input_valid),
    .io_iormac(bc_pe_796_io_iormac),
    .io_ve_out(bc_pe_796_io_ve_out),
    .io_ho_out(bc_pe_796_io_ho_out),
    .io_res_out(bc_pe_796_io_res_out)
  );
  bc_pe bc_pe_797 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_797_clock),
    .reset(bc_pe_797_reset),
    .io_ho_input(bc_pe_797_io_ho_input),
    .io_ve_input(bc_pe_797_io_ve_input),
    .io_input_valid(bc_pe_797_io_input_valid),
    .io_iormac(bc_pe_797_io_iormac),
    .io_ve_out(bc_pe_797_io_ve_out),
    .io_ho_out(bc_pe_797_io_ho_out),
    .io_res_out(bc_pe_797_io_res_out)
  );
  bc_pe bc_pe_798 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_798_clock),
    .reset(bc_pe_798_reset),
    .io_ho_input(bc_pe_798_io_ho_input),
    .io_ve_input(bc_pe_798_io_ve_input),
    .io_input_valid(bc_pe_798_io_input_valid),
    .io_iormac(bc_pe_798_io_iormac),
    .io_ve_out(bc_pe_798_io_ve_out),
    .io_ho_out(bc_pe_798_io_ho_out),
    .io_res_out(bc_pe_798_io_res_out)
  );
  bc_pe bc_pe_799 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_799_clock),
    .reset(bc_pe_799_reset),
    .io_ho_input(bc_pe_799_io_ho_input),
    .io_ve_input(bc_pe_799_io_ve_input),
    .io_input_valid(bc_pe_799_io_input_valid),
    .io_iormac(bc_pe_799_io_iormac),
    .io_ve_out(bc_pe_799_io_ve_out),
    .io_ho_out(bc_pe_799_io_ho_out),
    .io_res_out(bc_pe_799_io_res_out)
  );
  bc_pe bc_pe_800 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_800_clock),
    .reset(bc_pe_800_reset),
    .io_ho_input(bc_pe_800_io_ho_input),
    .io_ve_input(bc_pe_800_io_ve_input),
    .io_input_valid(bc_pe_800_io_input_valid),
    .io_iormac(bc_pe_800_io_iormac),
    .io_ve_out(bc_pe_800_io_ve_out),
    .io_ho_out(bc_pe_800_io_ho_out),
    .io_res_out(bc_pe_800_io_res_out)
  );
  bc_pe bc_pe_801 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_801_clock),
    .reset(bc_pe_801_reset),
    .io_ho_input(bc_pe_801_io_ho_input),
    .io_ve_input(bc_pe_801_io_ve_input),
    .io_input_valid(bc_pe_801_io_input_valid),
    .io_iormac(bc_pe_801_io_iormac),
    .io_ve_out(bc_pe_801_io_ve_out),
    .io_ho_out(bc_pe_801_io_ho_out),
    .io_res_out(bc_pe_801_io_res_out)
  );
  bc_pe bc_pe_802 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_802_clock),
    .reset(bc_pe_802_reset),
    .io_ho_input(bc_pe_802_io_ho_input),
    .io_ve_input(bc_pe_802_io_ve_input),
    .io_input_valid(bc_pe_802_io_input_valid),
    .io_iormac(bc_pe_802_io_iormac),
    .io_ve_out(bc_pe_802_io_ve_out),
    .io_ho_out(bc_pe_802_io_ho_out),
    .io_res_out(bc_pe_802_io_res_out)
  );
  bc_pe bc_pe_803 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_803_clock),
    .reset(bc_pe_803_reset),
    .io_ho_input(bc_pe_803_io_ho_input),
    .io_ve_input(bc_pe_803_io_ve_input),
    .io_input_valid(bc_pe_803_io_input_valid),
    .io_iormac(bc_pe_803_io_iormac),
    .io_ve_out(bc_pe_803_io_ve_out),
    .io_ho_out(bc_pe_803_io_ho_out),
    .io_res_out(bc_pe_803_io_res_out)
  );
  bc_pe bc_pe_804 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_804_clock),
    .reset(bc_pe_804_reset),
    .io_ho_input(bc_pe_804_io_ho_input),
    .io_ve_input(bc_pe_804_io_ve_input),
    .io_input_valid(bc_pe_804_io_input_valid),
    .io_iormac(bc_pe_804_io_iormac),
    .io_ve_out(bc_pe_804_io_ve_out),
    .io_ho_out(bc_pe_804_io_ho_out),
    .io_res_out(bc_pe_804_io_res_out)
  );
  bc_pe bc_pe_805 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_805_clock),
    .reset(bc_pe_805_reset),
    .io_ho_input(bc_pe_805_io_ho_input),
    .io_ve_input(bc_pe_805_io_ve_input),
    .io_input_valid(bc_pe_805_io_input_valid),
    .io_iormac(bc_pe_805_io_iormac),
    .io_ve_out(bc_pe_805_io_ve_out),
    .io_ho_out(bc_pe_805_io_ho_out),
    .io_res_out(bc_pe_805_io_res_out)
  );
  bc_pe bc_pe_806 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_806_clock),
    .reset(bc_pe_806_reset),
    .io_ho_input(bc_pe_806_io_ho_input),
    .io_ve_input(bc_pe_806_io_ve_input),
    .io_input_valid(bc_pe_806_io_input_valid),
    .io_iormac(bc_pe_806_io_iormac),
    .io_ve_out(bc_pe_806_io_ve_out),
    .io_ho_out(bc_pe_806_io_ho_out),
    .io_res_out(bc_pe_806_io_res_out)
  );
  bc_pe bc_pe_807 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_807_clock),
    .reset(bc_pe_807_reset),
    .io_ho_input(bc_pe_807_io_ho_input),
    .io_ve_input(bc_pe_807_io_ve_input),
    .io_input_valid(bc_pe_807_io_input_valid),
    .io_iormac(bc_pe_807_io_iormac),
    .io_ve_out(bc_pe_807_io_ve_out),
    .io_ho_out(bc_pe_807_io_ho_out),
    .io_res_out(bc_pe_807_io_res_out)
  );
  bc_pe bc_pe_808 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_808_clock),
    .reset(bc_pe_808_reset),
    .io_ho_input(bc_pe_808_io_ho_input),
    .io_ve_input(bc_pe_808_io_ve_input),
    .io_input_valid(bc_pe_808_io_input_valid),
    .io_iormac(bc_pe_808_io_iormac),
    .io_ve_out(bc_pe_808_io_ve_out),
    .io_ho_out(bc_pe_808_io_ho_out),
    .io_res_out(bc_pe_808_io_res_out)
  );
  bc_pe bc_pe_809 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_809_clock),
    .reset(bc_pe_809_reset),
    .io_ho_input(bc_pe_809_io_ho_input),
    .io_ve_input(bc_pe_809_io_ve_input),
    .io_input_valid(bc_pe_809_io_input_valid),
    .io_iormac(bc_pe_809_io_iormac),
    .io_ve_out(bc_pe_809_io_ve_out),
    .io_ho_out(bc_pe_809_io_ho_out),
    .io_res_out(bc_pe_809_io_res_out)
  );
  bc_pe bc_pe_810 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_810_clock),
    .reset(bc_pe_810_reset),
    .io_ho_input(bc_pe_810_io_ho_input),
    .io_ve_input(bc_pe_810_io_ve_input),
    .io_input_valid(bc_pe_810_io_input_valid),
    .io_iormac(bc_pe_810_io_iormac),
    .io_ve_out(bc_pe_810_io_ve_out),
    .io_ho_out(bc_pe_810_io_ho_out),
    .io_res_out(bc_pe_810_io_res_out)
  );
  bc_pe bc_pe_811 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_811_clock),
    .reset(bc_pe_811_reset),
    .io_ho_input(bc_pe_811_io_ho_input),
    .io_ve_input(bc_pe_811_io_ve_input),
    .io_input_valid(bc_pe_811_io_input_valid),
    .io_iormac(bc_pe_811_io_iormac),
    .io_ve_out(bc_pe_811_io_ve_out),
    .io_ho_out(bc_pe_811_io_ho_out),
    .io_res_out(bc_pe_811_io_res_out)
  );
  bc_pe bc_pe_812 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_812_clock),
    .reset(bc_pe_812_reset),
    .io_ho_input(bc_pe_812_io_ho_input),
    .io_ve_input(bc_pe_812_io_ve_input),
    .io_input_valid(bc_pe_812_io_input_valid),
    .io_iormac(bc_pe_812_io_iormac),
    .io_ve_out(bc_pe_812_io_ve_out),
    .io_ho_out(bc_pe_812_io_ho_out),
    .io_res_out(bc_pe_812_io_res_out)
  );
  bc_pe bc_pe_813 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_813_clock),
    .reset(bc_pe_813_reset),
    .io_ho_input(bc_pe_813_io_ho_input),
    .io_ve_input(bc_pe_813_io_ve_input),
    .io_input_valid(bc_pe_813_io_input_valid),
    .io_iormac(bc_pe_813_io_iormac),
    .io_ve_out(bc_pe_813_io_ve_out),
    .io_ho_out(bc_pe_813_io_ho_out),
    .io_res_out(bc_pe_813_io_res_out)
  );
  bc_pe bc_pe_814 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_814_clock),
    .reset(bc_pe_814_reset),
    .io_ho_input(bc_pe_814_io_ho_input),
    .io_ve_input(bc_pe_814_io_ve_input),
    .io_input_valid(bc_pe_814_io_input_valid),
    .io_iormac(bc_pe_814_io_iormac),
    .io_ve_out(bc_pe_814_io_ve_out),
    .io_ho_out(bc_pe_814_io_ho_out),
    .io_res_out(bc_pe_814_io_res_out)
  );
  bc_pe bc_pe_815 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_815_clock),
    .reset(bc_pe_815_reset),
    .io_ho_input(bc_pe_815_io_ho_input),
    .io_ve_input(bc_pe_815_io_ve_input),
    .io_input_valid(bc_pe_815_io_input_valid),
    .io_iormac(bc_pe_815_io_iormac),
    .io_ve_out(bc_pe_815_io_ve_out),
    .io_ho_out(bc_pe_815_io_ho_out),
    .io_res_out(bc_pe_815_io_res_out)
  );
  bc_pe bc_pe_816 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_816_clock),
    .reset(bc_pe_816_reset),
    .io_ho_input(bc_pe_816_io_ho_input),
    .io_ve_input(bc_pe_816_io_ve_input),
    .io_input_valid(bc_pe_816_io_input_valid),
    .io_iormac(bc_pe_816_io_iormac),
    .io_ve_out(bc_pe_816_io_ve_out),
    .io_ho_out(bc_pe_816_io_ho_out),
    .io_res_out(bc_pe_816_io_res_out)
  );
  bc_pe bc_pe_817 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_817_clock),
    .reset(bc_pe_817_reset),
    .io_ho_input(bc_pe_817_io_ho_input),
    .io_ve_input(bc_pe_817_io_ve_input),
    .io_input_valid(bc_pe_817_io_input_valid),
    .io_iormac(bc_pe_817_io_iormac),
    .io_ve_out(bc_pe_817_io_ve_out),
    .io_ho_out(bc_pe_817_io_ho_out),
    .io_res_out(bc_pe_817_io_res_out)
  );
  bc_pe bc_pe_818 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_818_clock),
    .reset(bc_pe_818_reset),
    .io_ho_input(bc_pe_818_io_ho_input),
    .io_ve_input(bc_pe_818_io_ve_input),
    .io_input_valid(bc_pe_818_io_input_valid),
    .io_iormac(bc_pe_818_io_iormac),
    .io_ve_out(bc_pe_818_io_ve_out),
    .io_ho_out(bc_pe_818_io_ho_out),
    .io_res_out(bc_pe_818_io_res_out)
  );
  bc_pe bc_pe_819 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_819_clock),
    .reset(bc_pe_819_reset),
    .io_ho_input(bc_pe_819_io_ho_input),
    .io_ve_input(bc_pe_819_io_ve_input),
    .io_input_valid(bc_pe_819_io_input_valid),
    .io_iormac(bc_pe_819_io_iormac),
    .io_ve_out(bc_pe_819_io_ve_out),
    .io_ho_out(bc_pe_819_io_ho_out),
    .io_res_out(bc_pe_819_io_res_out)
  );
  bc_pe bc_pe_820 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_820_clock),
    .reset(bc_pe_820_reset),
    .io_ho_input(bc_pe_820_io_ho_input),
    .io_ve_input(bc_pe_820_io_ve_input),
    .io_input_valid(bc_pe_820_io_input_valid),
    .io_iormac(bc_pe_820_io_iormac),
    .io_ve_out(bc_pe_820_io_ve_out),
    .io_ho_out(bc_pe_820_io_ho_out),
    .io_res_out(bc_pe_820_io_res_out)
  );
  bc_pe bc_pe_821 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_821_clock),
    .reset(bc_pe_821_reset),
    .io_ho_input(bc_pe_821_io_ho_input),
    .io_ve_input(bc_pe_821_io_ve_input),
    .io_input_valid(bc_pe_821_io_input_valid),
    .io_iormac(bc_pe_821_io_iormac),
    .io_ve_out(bc_pe_821_io_ve_out),
    .io_ho_out(bc_pe_821_io_ho_out),
    .io_res_out(bc_pe_821_io_res_out)
  );
  bc_pe bc_pe_822 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_822_clock),
    .reset(bc_pe_822_reset),
    .io_ho_input(bc_pe_822_io_ho_input),
    .io_ve_input(bc_pe_822_io_ve_input),
    .io_input_valid(bc_pe_822_io_input_valid),
    .io_iormac(bc_pe_822_io_iormac),
    .io_ve_out(bc_pe_822_io_ve_out),
    .io_ho_out(bc_pe_822_io_ho_out),
    .io_res_out(bc_pe_822_io_res_out)
  );
  bc_pe bc_pe_823 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_823_clock),
    .reset(bc_pe_823_reset),
    .io_ho_input(bc_pe_823_io_ho_input),
    .io_ve_input(bc_pe_823_io_ve_input),
    .io_input_valid(bc_pe_823_io_input_valid),
    .io_iormac(bc_pe_823_io_iormac),
    .io_ve_out(bc_pe_823_io_ve_out),
    .io_ho_out(bc_pe_823_io_ho_out),
    .io_res_out(bc_pe_823_io_res_out)
  );
  bc_pe bc_pe_824 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_824_clock),
    .reset(bc_pe_824_reset),
    .io_ho_input(bc_pe_824_io_ho_input),
    .io_ve_input(bc_pe_824_io_ve_input),
    .io_input_valid(bc_pe_824_io_input_valid),
    .io_iormac(bc_pe_824_io_iormac),
    .io_ve_out(bc_pe_824_io_ve_out),
    .io_ho_out(bc_pe_824_io_ho_out),
    .io_res_out(bc_pe_824_io_res_out)
  );
  bc_pe bc_pe_825 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_825_clock),
    .reset(bc_pe_825_reset),
    .io_ho_input(bc_pe_825_io_ho_input),
    .io_ve_input(bc_pe_825_io_ve_input),
    .io_input_valid(bc_pe_825_io_input_valid),
    .io_iormac(bc_pe_825_io_iormac),
    .io_ve_out(bc_pe_825_io_ve_out),
    .io_ho_out(bc_pe_825_io_ho_out),
    .io_res_out(bc_pe_825_io_res_out)
  );
  bc_pe bc_pe_826 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_826_clock),
    .reset(bc_pe_826_reset),
    .io_ho_input(bc_pe_826_io_ho_input),
    .io_ve_input(bc_pe_826_io_ve_input),
    .io_input_valid(bc_pe_826_io_input_valid),
    .io_iormac(bc_pe_826_io_iormac),
    .io_ve_out(bc_pe_826_io_ve_out),
    .io_ho_out(bc_pe_826_io_ho_out),
    .io_res_out(bc_pe_826_io_res_out)
  );
  bc_pe bc_pe_827 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_827_clock),
    .reset(bc_pe_827_reset),
    .io_ho_input(bc_pe_827_io_ho_input),
    .io_ve_input(bc_pe_827_io_ve_input),
    .io_input_valid(bc_pe_827_io_input_valid),
    .io_iormac(bc_pe_827_io_iormac),
    .io_ve_out(bc_pe_827_io_ve_out),
    .io_ho_out(bc_pe_827_io_ho_out),
    .io_res_out(bc_pe_827_io_res_out)
  );
  bc_pe bc_pe_828 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_828_clock),
    .reset(bc_pe_828_reset),
    .io_ho_input(bc_pe_828_io_ho_input),
    .io_ve_input(bc_pe_828_io_ve_input),
    .io_input_valid(bc_pe_828_io_input_valid),
    .io_iormac(bc_pe_828_io_iormac),
    .io_ve_out(bc_pe_828_io_ve_out),
    .io_ho_out(bc_pe_828_io_ho_out),
    .io_res_out(bc_pe_828_io_res_out)
  );
  bc_pe bc_pe_829 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_829_clock),
    .reset(bc_pe_829_reset),
    .io_ho_input(bc_pe_829_io_ho_input),
    .io_ve_input(bc_pe_829_io_ve_input),
    .io_input_valid(bc_pe_829_io_input_valid),
    .io_iormac(bc_pe_829_io_iormac),
    .io_ve_out(bc_pe_829_io_ve_out),
    .io_ho_out(bc_pe_829_io_ho_out),
    .io_res_out(bc_pe_829_io_res_out)
  );
  bc_pe bc_pe_830 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_830_clock),
    .reset(bc_pe_830_reset),
    .io_ho_input(bc_pe_830_io_ho_input),
    .io_ve_input(bc_pe_830_io_ve_input),
    .io_input_valid(bc_pe_830_io_input_valid),
    .io_iormac(bc_pe_830_io_iormac),
    .io_ve_out(bc_pe_830_io_ve_out),
    .io_ho_out(bc_pe_830_io_ho_out),
    .io_res_out(bc_pe_830_io_res_out)
  );
  bc_pe bc_pe_831 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_831_clock),
    .reset(bc_pe_831_reset),
    .io_ho_input(bc_pe_831_io_ho_input),
    .io_ve_input(bc_pe_831_io_ve_input),
    .io_input_valid(bc_pe_831_io_input_valid),
    .io_iormac(bc_pe_831_io_iormac),
    .io_ve_out(bc_pe_831_io_ve_out),
    .io_ho_out(bc_pe_831_io_ho_out),
    .io_res_out(bc_pe_831_io_res_out)
  );
  bc_pe bc_pe_832 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_832_clock),
    .reset(bc_pe_832_reset),
    .io_ho_input(bc_pe_832_io_ho_input),
    .io_ve_input(bc_pe_832_io_ve_input),
    .io_input_valid(bc_pe_832_io_input_valid),
    .io_iormac(bc_pe_832_io_iormac),
    .io_ve_out(bc_pe_832_io_ve_out),
    .io_ho_out(bc_pe_832_io_ho_out),
    .io_res_out(bc_pe_832_io_res_out)
  );
  bc_pe bc_pe_833 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_833_clock),
    .reset(bc_pe_833_reset),
    .io_ho_input(bc_pe_833_io_ho_input),
    .io_ve_input(bc_pe_833_io_ve_input),
    .io_input_valid(bc_pe_833_io_input_valid),
    .io_iormac(bc_pe_833_io_iormac),
    .io_ve_out(bc_pe_833_io_ve_out),
    .io_ho_out(bc_pe_833_io_ho_out),
    .io_res_out(bc_pe_833_io_res_out)
  );
  bc_pe bc_pe_834 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_834_clock),
    .reset(bc_pe_834_reset),
    .io_ho_input(bc_pe_834_io_ho_input),
    .io_ve_input(bc_pe_834_io_ve_input),
    .io_input_valid(bc_pe_834_io_input_valid),
    .io_iormac(bc_pe_834_io_iormac),
    .io_ve_out(bc_pe_834_io_ve_out),
    .io_ho_out(bc_pe_834_io_ho_out),
    .io_res_out(bc_pe_834_io_res_out)
  );
  bc_pe bc_pe_835 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_835_clock),
    .reset(bc_pe_835_reset),
    .io_ho_input(bc_pe_835_io_ho_input),
    .io_ve_input(bc_pe_835_io_ve_input),
    .io_input_valid(bc_pe_835_io_input_valid),
    .io_iormac(bc_pe_835_io_iormac),
    .io_ve_out(bc_pe_835_io_ve_out),
    .io_ho_out(bc_pe_835_io_ho_out),
    .io_res_out(bc_pe_835_io_res_out)
  );
  bc_pe bc_pe_836 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_836_clock),
    .reset(bc_pe_836_reset),
    .io_ho_input(bc_pe_836_io_ho_input),
    .io_ve_input(bc_pe_836_io_ve_input),
    .io_input_valid(bc_pe_836_io_input_valid),
    .io_iormac(bc_pe_836_io_iormac),
    .io_ve_out(bc_pe_836_io_ve_out),
    .io_ho_out(bc_pe_836_io_ho_out),
    .io_res_out(bc_pe_836_io_res_out)
  );
  bc_pe bc_pe_837 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_837_clock),
    .reset(bc_pe_837_reset),
    .io_ho_input(bc_pe_837_io_ho_input),
    .io_ve_input(bc_pe_837_io_ve_input),
    .io_input_valid(bc_pe_837_io_input_valid),
    .io_iormac(bc_pe_837_io_iormac),
    .io_ve_out(bc_pe_837_io_ve_out),
    .io_ho_out(bc_pe_837_io_ho_out),
    .io_res_out(bc_pe_837_io_res_out)
  );
  bc_pe bc_pe_838 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_838_clock),
    .reset(bc_pe_838_reset),
    .io_ho_input(bc_pe_838_io_ho_input),
    .io_ve_input(bc_pe_838_io_ve_input),
    .io_input_valid(bc_pe_838_io_input_valid),
    .io_iormac(bc_pe_838_io_iormac),
    .io_ve_out(bc_pe_838_io_ve_out),
    .io_ho_out(bc_pe_838_io_ho_out),
    .io_res_out(bc_pe_838_io_res_out)
  );
  bc_pe bc_pe_839 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_839_clock),
    .reset(bc_pe_839_reset),
    .io_ho_input(bc_pe_839_io_ho_input),
    .io_ve_input(bc_pe_839_io_ve_input),
    .io_input_valid(bc_pe_839_io_input_valid),
    .io_iormac(bc_pe_839_io_iormac),
    .io_ve_out(bc_pe_839_io_ve_out),
    .io_ho_out(bc_pe_839_io_ho_out),
    .io_res_out(bc_pe_839_io_res_out)
  );
  bc_pe bc_pe_840 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_840_clock),
    .reset(bc_pe_840_reset),
    .io_ho_input(bc_pe_840_io_ho_input),
    .io_ve_input(bc_pe_840_io_ve_input),
    .io_input_valid(bc_pe_840_io_input_valid),
    .io_iormac(bc_pe_840_io_iormac),
    .io_ve_out(bc_pe_840_io_ve_out),
    .io_ho_out(bc_pe_840_io_ho_out),
    .io_res_out(bc_pe_840_io_res_out)
  );
  bc_pe bc_pe_841 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_841_clock),
    .reset(bc_pe_841_reset),
    .io_ho_input(bc_pe_841_io_ho_input),
    .io_ve_input(bc_pe_841_io_ve_input),
    .io_input_valid(bc_pe_841_io_input_valid),
    .io_iormac(bc_pe_841_io_iormac),
    .io_ve_out(bc_pe_841_io_ve_out),
    .io_ho_out(bc_pe_841_io_ho_out),
    .io_res_out(bc_pe_841_io_res_out)
  );
  bc_pe bc_pe_842 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_842_clock),
    .reset(bc_pe_842_reset),
    .io_ho_input(bc_pe_842_io_ho_input),
    .io_ve_input(bc_pe_842_io_ve_input),
    .io_input_valid(bc_pe_842_io_input_valid),
    .io_iormac(bc_pe_842_io_iormac),
    .io_ve_out(bc_pe_842_io_ve_out),
    .io_ho_out(bc_pe_842_io_ho_out),
    .io_res_out(bc_pe_842_io_res_out)
  );
  bc_pe bc_pe_843 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_843_clock),
    .reset(bc_pe_843_reset),
    .io_ho_input(bc_pe_843_io_ho_input),
    .io_ve_input(bc_pe_843_io_ve_input),
    .io_input_valid(bc_pe_843_io_input_valid),
    .io_iormac(bc_pe_843_io_iormac),
    .io_ve_out(bc_pe_843_io_ve_out),
    .io_ho_out(bc_pe_843_io_ho_out),
    .io_res_out(bc_pe_843_io_res_out)
  );
  bc_pe bc_pe_844 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_844_clock),
    .reset(bc_pe_844_reset),
    .io_ho_input(bc_pe_844_io_ho_input),
    .io_ve_input(bc_pe_844_io_ve_input),
    .io_input_valid(bc_pe_844_io_input_valid),
    .io_iormac(bc_pe_844_io_iormac),
    .io_ve_out(bc_pe_844_io_ve_out),
    .io_ho_out(bc_pe_844_io_ho_out),
    .io_res_out(bc_pe_844_io_res_out)
  );
  bc_pe bc_pe_845 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_845_clock),
    .reset(bc_pe_845_reset),
    .io_ho_input(bc_pe_845_io_ho_input),
    .io_ve_input(bc_pe_845_io_ve_input),
    .io_input_valid(bc_pe_845_io_input_valid),
    .io_iormac(bc_pe_845_io_iormac),
    .io_ve_out(bc_pe_845_io_ve_out),
    .io_ho_out(bc_pe_845_io_ho_out),
    .io_res_out(bc_pe_845_io_res_out)
  );
  bc_pe bc_pe_846 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_846_clock),
    .reset(bc_pe_846_reset),
    .io_ho_input(bc_pe_846_io_ho_input),
    .io_ve_input(bc_pe_846_io_ve_input),
    .io_input_valid(bc_pe_846_io_input_valid),
    .io_iormac(bc_pe_846_io_iormac),
    .io_ve_out(bc_pe_846_io_ve_out),
    .io_ho_out(bc_pe_846_io_ho_out),
    .io_res_out(bc_pe_846_io_res_out)
  );
  bc_pe bc_pe_847 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_847_clock),
    .reset(bc_pe_847_reset),
    .io_ho_input(bc_pe_847_io_ho_input),
    .io_ve_input(bc_pe_847_io_ve_input),
    .io_input_valid(bc_pe_847_io_input_valid),
    .io_iormac(bc_pe_847_io_iormac),
    .io_ve_out(bc_pe_847_io_ve_out),
    .io_ho_out(bc_pe_847_io_ho_out),
    .io_res_out(bc_pe_847_io_res_out)
  );
  bc_pe bc_pe_848 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_848_clock),
    .reset(bc_pe_848_reset),
    .io_ho_input(bc_pe_848_io_ho_input),
    .io_ve_input(bc_pe_848_io_ve_input),
    .io_input_valid(bc_pe_848_io_input_valid),
    .io_iormac(bc_pe_848_io_iormac),
    .io_ve_out(bc_pe_848_io_ve_out),
    .io_ho_out(bc_pe_848_io_ho_out),
    .io_res_out(bc_pe_848_io_res_out)
  );
  bc_pe bc_pe_849 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_849_clock),
    .reset(bc_pe_849_reset),
    .io_ho_input(bc_pe_849_io_ho_input),
    .io_ve_input(bc_pe_849_io_ve_input),
    .io_input_valid(bc_pe_849_io_input_valid),
    .io_iormac(bc_pe_849_io_iormac),
    .io_ve_out(bc_pe_849_io_ve_out),
    .io_ho_out(bc_pe_849_io_ho_out),
    .io_res_out(bc_pe_849_io_res_out)
  );
  bc_pe bc_pe_850 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_850_clock),
    .reset(bc_pe_850_reset),
    .io_ho_input(bc_pe_850_io_ho_input),
    .io_ve_input(bc_pe_850_io_ve_input),
    .io_input_valid(bc_pe_850_io_input_valid),
    .io_iormac(bc_pe_850_io_iormac),
    .io_ve_out(bc_pe_850_io_ve_out),
    .io_ho_out(bc_pe_850_io_ho_out),
    .io_res_out(bc_pe_850_io_res_out)
  );
  bc_pe bc_pe_851 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_851_clock),
    .reset(bc_pe_851_reset),
    .io_ho_input(bc_pe_851_io_ho_input),
    .io_ve_input(bc_pe_851_io_ve_input),
    .io_input_valid(bc_pe_851_io_input_valid),
    .io_iormac(bc_pe_851_io_iormac),
    .io_ve_out(bc_pe_851_io_ve_out),
    .io_ho_out(bc_pe_851_io_ho_out),
    .io_res_out(bc_pe_851_io_res_out)
  );
  bc_pe bc_pe_852 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_852_clock),
    .reset(bc_pe_852_reset),
    .io_ho_input(bc_pe_852_io_ho_input),
    .io_ve_input(bc_pe_852_io_ve_input),
    .io_input_valid(bc_pe_852_io_input_valid),
    .io_iormac(bc_pe_852_io_iormac),
    .io_ve_out(bc_pe_852_io_ve_out),
    .io_ho_out(bc_pe_852_io_ho_out),
    .io_res_out(bc_pe_852_io_res_out)
  );
  bc_pe bc_pe_853 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_853_clock),
    .reset(bc_pe_853_reset),
    .io_ho_input(bc_pe_853_io_ho_input),
    .io_ve_input(bc_pe_853_io_ve_input),
    .io_input_valid(bc_pe_853_io_input_valid),
    .io_iormac(bc_pe_853_io_iormac),
    .io_ve_out(bc_pe_853_io_ve_out),
    .io_ho_out(bc_pe_853_io_ho_out),
    .io_res_out(bc_pe_853_io_res_out)
  );
  bc_pe bc_pe_854 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_854_clock),
    .reset(bc_pe_854_reset),
    .io_ho_input(bc_pe_854_io_ho_input),
    .io_ve_input(bc_pe_854_io_ve_input),
    .io_input_valid(bc_pe_854_io_input_valid),
    .io_iormac(bc_pe_854_io_iormac),
    .io_ve_out(bc_pe_854_io_ve_out),
    .io_ho_out(bc_pe_854_io_ho_out),
    .io_res_out(bc_pe_854_io_res_out)
  );
  bc_pe bc_pe_855 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_855_clock),
    .reset(bc_pe_855_reset),
    .io_ho_input(bc_pe_855_io_ho_input),
    .io_ve_input(bc_pe_855_io_ve_input),
    .io_input_valid(bc_pe_855_io_input_valid),
    .io_iormac(bc_pe_855_io_iormac),
    .io_ve_out(bc_pe_855_io_ve_out),
    .io_ho_out(bc_pe_855_io_ho_out),
    .io_res_out(bc_pe_855_io_res_out)
  );
  bc_pe bc_pe_856 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_856_clock),
    .reset(bc_pe_856_reset),
    .io_ho_input(bc_pe_856_io_ho_input),
    .io_ve_input(bc_pe_856_io_ve_input),
    .io_input_valid(bc_pe_856_io_input_valid),
    .io_iormac(bc_pe_856_io_iormac),
    .io_ve_out(bc_pe_856_io_ve_out),
    .io_ho_out(bc_pe_856_io_ho_out),
    .io_res_out(bc_pe_856_io_res_out)
  );
  bc_pe bc_pe_857 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_857_clock),
    .reset(bc_pe_857_reset),
    .io_ho_input(bc_pe_857_io_ho_input),
    .io_ve_input(bc_pe_857_io_ve_input),
    .io_input_valid(bc_pe_857_io_input_valid),
    .io_iormac(bc_pe_857_io_iormac),
    .io_ve_out(bc_pe_857_io_ve_out),
    .io_ho_out(bc_pe_857_io_ho_out),
    .io_res_out(bc_pe_857_io_res_out)
  );
  bc_pe bc_pe_858 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_858_clock),
    .reset(bc_pe_858_reset),
    .io_ho_input(bc_pe_858_io_ho_input),
    .io_ve_input(bc_pe_858_io_ve_input),
    .io_input_valid(bc_pe_858_io_input_valid),
    .io_iormac(bc_pe_858_io_iormac),
    .io_ve_out(bc_pe_858_io_ve_out),
    .io_ho_out(bc_pe_858_io_ho_out),
    .io_res_out(bc_pe_858_io_res_out)
  );
  bc_pe bc_pe_859 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_859_clock),
    .reset(bc_pe_859_reset),
    .io_ho_input(bc_pe_859_io_ho_input),
    .io_ve_input(bc_pe_859_io_ve_input),
    .io_input_valid(bc_pe_859_io_input_valid),
    .io_iormac(bc_pe_859_io_iormac),
    .io_ve_out(bc_pe_859_io_ve_out),
    .io_ho_out(bc_pe_859_io_ho_out),
    .io_res_out(bc_pe_859_io_res_out)
  );
  bc_pe bc_pe_860 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_860_clock),
    .reset(bc_pe_860_reset),
    .io_ho_input(bc_pe_860_io_ho_input),
    .io_ve_input(bc_pe_860_io_ve_input),
    .io_input_valid(bc_pe_860_io_input_valid),
    .io_iormac(bc_pe_860_io_iormac),
    .io_ve_out(bc_pe_860_io_ve_out),
    .io_ho_out(bc_pe_860_io_ho_out),
    .io_res_out(bc_pe_860_io_res_out)
  );
  bc_pe bc_pe_861 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_861_clock),
    .reset(bc_pe_861_reset),
    .io_ho_input(bc_pe_861_io_ho_input),
    .io_ve_input(bc_pe_861_io_ve_input),
    .io_input_valid(bc_pe_861_io_input_valid),
    .io_iormac(bc_pe_861_io_iormac),
    .io_ve_out(bc_pe_861_io_ve_out),
    .io_ho_out(bc_pe_861_io_ho_out),
    .io_res_out(bc_pe_861_io_res_out)
  );
  bc_pe bc_pe_862 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_862_clock),
    .reset(bc_pe_862_reset),
    .io_ho_input(bc_pe_862_io_ho_input),
    .io_ve_input(bc_pe_862_io_ve_input),
    .io_input_valid(bc_pe_862_io_input_valid),
    .io_iormac(bc_pe_862_io_iormac),
    .io_ve_out(bc_pe_862_io_ve_out),
    .io_ho_out(bc_pe_862_io_ho_out),
    .io_res_out(bc_pe_862_io_res_out)
  );
  bc_pe bc_pe_863 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_863_clock),
    .reset(bc_pe_863_reset),
    .io_ho_input(bc_pe_863_io_ho_input),
    .io_ve_input(bc_pe_863_io_ve_input),
    .io_input_valid(bc_pe_863_io_input_valid),
    .io_iormac(bc_pe_863_io_iormac),
    .io_ve_out(bc_pe_863_io_ve_out),
    .io_ho_out(bc_pe_863_io_ho_out),
    .io_res_out(bc_pe_863_io_res_out)
  );
  bc_pe bc_pe_864 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_864_clock),
    .reset(bc_pe_864_reset),
    .io_ho_input(bc_pe_864_io_ho_input),
    .io_ve_input(bc_pe_864_io_ve_input),
    .io_input_valid(bc_pe_864_io_input_valid),
    .io_iormac(bc_pe_864_io_iormac),
    .io_ve_out(bc_pe_864_io_ve_out),
    .io_ho_out(bc_pe_864_io_ho_out),
    .io_res_out(bc_pe_864_io_res_out)
  );
  bc_pe bc_pe_865 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_865_clock),
    .reset(bc_pe_865_reset),
    .io_ho_input(bc_pe_865_io_ho_input),
    .io_ve_input(bc_pe_865_io_ve_input),
    .io_input_valid(bc_pe_865_io_input_valid),
    .io_iormac(bc_pe_865_io_iormac),
    .io_ve_out(bc_pe_865_io_ve_out),
    .io_ho_out(bc_pe_865_io_ho_out),
    .io_res_out(bc_pe_865_io_res_out)
  );
  bc_pe bc_pe_866 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_866_clock),
    .reset(bc_pe_866_reset),
    .io_ho_input(bc_pe_866_io_ho_input),
    .io_ve_input(bc_pe_866_io_ve_input),
    .io_input_valid(bc_pe_866_io_input_valid),
    .io_iormac(bc_pe_866_io_iormac),
    .io_ve_out(bc_pe_866_io_ve_out),
    .io_ho_out(bc_pe_866_io_ho_out),
    .io_res_out(bc_pe_866_io_res_out)
  );
  bc_pe bc_pe_867 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_867_clock),
    .reset(bc_pe_867_reset),
    .io_ho_input(bc_pe_867_io_ho_input),
    .io_ve_input(bc_pe_867_io_ve_input),
    .io_input_valid(bc_pe_867_io_input_valid),
    .io_iormac(bc_pe_867_io_iormac),
    .io_ve_out(bc_pe_867_io_ve_out),
    .io_ho_out(bc_pe_867_io_ho_out),
    .io_res_out(bc_pe_867_io_res_out)
  );
  bc_pe bc_pe_868 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_868_clock),
    .reset(bc_pe_868_reset),
    .io_ho_input(bc_pe_868_io_ho_input),
    .io_ve_input(bc_pe_868_io_ve_input),
    .io_input_valid(bc_pe_868_io_input_valid),
    .io_iormac(bc_pe_868_io_iormac),
    .io_ve_out(bc_pe_868_io_ve_out),
    .io_ho_out(bc_pe_868_io_ho_out),
    .io_res_out(bc_pe_868_io_res_out)
  );
  bc_pe bc_pe_869 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_869_clock),
    .reset(bc_pe_869_reset),
    .io_ho_input(bc_pe_869_io_ho_input),
    .io_ve_input(bc_pe_869_io_ve_input),
    .io_input_valid(bc_pe_869_io_input_valid),
    .io_iormac(bc_pe_869_io_iormac),
    .io_ve_out(bc_pe_869_io_ve_out),
    .io_ho_out(bc_pe_869_io_ho_out),
    .io_res_out(bc_pe_869_io_res_out)
  );
  bc_pe bc_pe_870 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_870_clock),
    .reset(bc_pe_870_reset),
    .io_ho_input(bc_pe_870_io_ho_input),
    .io_ve_input(bc_pe_870_io_ve_input),
    .io_input_valid(bc_pe_870_io_input_valid),
    .io_iormac(bc_pe_870_io_iormac),
    .io_ve_out(bc_pe_870_io_ve_out),
    .io_ho_out(bc_pe_870_io_ho_out),
    .io_res_out(bc_pe_870_io_res_out)
  );
  bc_pe bc_pe_871 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_871_clock),
    .reset(bc_pe_871_reset),
    .io_ho_input(bc_pe_871_io_ho_input),
    .io_ve_input(bc_pe_871_io_ve_input),
    .io_input_valid(bc_pe_871_io_input_valid),
    .io_iormac(bc_pe_871_io_iormac),
    .io_ve_out(bc_pe_871_io_ve_out),
    .io_ho_out(bc_pe_871_io_ho_out),
    .io_res_out(bc_pe_871_io_res_out)
  );
  bc_pe bc_pe_872 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_872_clock),
    .reset(bc_pe_872_reset),
    .io_ho_input(bc_pe_872_io_ho_input),
    .io_ve_input(bc_pe_872_io_ve_input),
    .io_input_valid(bc_pe_872_io_input_valid),
    .io_iormac(bc_pe_872_io_iormac),
    .io_ve_out(bc_pe_872_io_ve_out),
    .io_ho_out(bc_pe_872_io_ho_out),
    .io_res_out(bc_pe_872_io_res_out)
  );
  bc_pe bc_pe_873 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_873_clock),
    .reset(bc_pe_873_reset),
    .io_ho_input(bc_pe_873_io_ho_input),
    .io_ve_input(bc_pe_873_io_ve_input),
    .io_input_valid(bc_pe_873_io_input_valid),
    .io_iormac(bc_pe_873_io_iormac),
    .io_ve_out(bc_pe_873_io_ve_out),
    .io_ho_out(bc_pe_873_io_ho_out),
    .io_res_out(bc_pe_873_io_res_out)
  );
  bc_pe bc_pe_874 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_874_clock),
    .reset(bc_pe_874_reset),
    .io_ho_input(bc_pe_874_io_ho_input),
    .io_ve_input(bc_pe_874_io_ve_input),
    .io_input_valid(bc_pe_874_io_input_valid),
    .io_iormac(bc_pe_874_io_iormac),
    .io_ve_out(bc_pe_874_io_ve_out),
    .io_ho_out(bc_pe_874_io_ho_out),
    .io_res_out(bc_pe_874_io_res_out)
  );
  bc_pe bc_pe_875 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_875_clock),
    .reset(bc_pe_875_reset),
    .io_ho_input(bc_pe_875_io_ho_input),
    .io_ve_input(bc_pe_875_io_ve_input),
    .io_input_valid(bc_pe_875_io_input_valid),
    .io_iormac(bc_pe_875_io_iormac),
    .io_ve_out(bc_pe_875_io_ve_out),
    .io_ho_out(bc_pe_875_io_ho_out),
    .io_res_out(bc_pe_875_io_res_out)
  );
  bc_pe bc_pe_876 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_876_clock),
    .reset(bc_pe_876_reset),
    .io_ho_input(bc_pe_876_io_ho_input),
    .io_ve_input(bc_pe_876_io_ve_input),
    .io_input_valid(bc_pe_876_io_input_valid),
    .io_iormac(bc_pe_876_io_iormac),
    .io_ve_out(bc_pe_876_io_ve_out),
    .io_ho_out(bc_pe_876_io_ho_out),
    .io_res_out(bc_pe_876_io_res_out)
  );
  bc_pe bc_pe_877 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_877_clock),
    .reset(bc_pe_877_reset),
    .io_ho_input(bc_pe_877_io_ho_input),
    .io_ve_input(bc_pe_877_io_ve_input),
    .io_input_valid(bc_pe_877_io_input_valid),
    .io_iormac(bc_pe_877_io_iormac),
    .io_ve_out(bc_pe_877_io_ve_out),
    .io_ho_out(bc_pe_877_io_ho_out),
    .io_res_out(bc_pe_877_io_res_out)
  );
  bc_pe bc_pe_878 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_878_clock),
    .reset(bc_pe_878_reset),
    .io_ho_input(bc_pe_878_io_ho_input),
    .io_ve_input(bc_pe_878_io_ve_input),
    .io_input_valid(bc_pe_878_io_input_valid),
    .io_iormac(bc_pe_878_io_iormac),
    .io_ve_out(bc_pe_878_io_ve_out),
    .io_ho_out(bc_pe_878_io_ho_out),
    .io_res_out(bc_pe_878_io_res_out)
  );
  bc_pe bc_pe_879 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_879_clock),
    .reset(bc_pe_879_reset),
    .io_ho_input(bc_pe_879_io_ho_input),
    .io_ve_input(bc_pe_879_io_ve_input),
    .io_input_valid(bc_pe_879_io_input_valid),
    .io_iormac(bc_pe_879_io_iormac),
    .io_ve_out(bc_pe_879_io_ve_out),
    .io_ho_out(bc_pe_879_io_ho_out),
    .io_res_out(bc_pe_879_io_res_out)
  );
  bc_pe bc_pe_880 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_880_clock),
    .reset(bc_pe_880_reset),
    .io_ho_input(bc_pe_880_io_ho_input),
    .io_ve_input(bc_pe_880_io_ve_input),
    .io_input_valid(bc_pe_880_io_input_valid),
    .io_iormac(bc_pe_880_io_iormac),
    .io_ve_out(bc_pe_880_io_ve_out),
    .io_ho_out(bc_pe_880_io_ho_out),
    .io_res_out(bc_pe_880_io_res_out)
  );
  bc_pe bc_pe_881 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_881_clock),
    .reset(bc_pe_881_reset),
    .io_ho_input(bc_pe_881_io_ho_input),
    .io_ve_input(bc_pe_881_io_ve_input),
    .io_input_valid(bc_pe_881_io_input_valid),
    .io_iormac(bc_pe_881_io_iormac),
    .io_ve_out(bc_pe_881_io_ve_out),
    .io_ho_out(bc_pe_881_io_ho_out),
    .io_res_out(bc_pe_881_io_res_out)
  );
  bc_pe bc_pe_882 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_882_clock),
    .reset(bc_pe_882_reset),
    .io_ho_input(bc_pe_882_io_ho_input),
    .io_ve_input(bc_pe_882_io_ve_input),
    .io_input_valid(bc_pe_882_io_input_valid),
    .io_iormac(bc_pe_882_io_iormac),
    .io_ve_out(bc_pe_882_io_ve_out),
    .io_ho_out(bc_pe_882_io_ho_out),
    .io_res_out(bc_pe_882_io_res_out)
  );
  bc_pe bc_pe_883 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_883_clock),
    .reset(bc_pe_883_reset),
    .io_ho_input(bc_pe_883_io_ho_input),
    .io_ve_input(bc_pe_883_io_ve_input),
    .io_input_valid(bc_pe_883_io_input_valid),
    .io_iormac(bc_pe_883_io_iormac),
    .io_ve_out(bc_pe_883_io_ve_out),
    .io_ho_out(bc_pe_883_io_ho_out),
    .io_res_out(bc_pe_883_io_res_out)
  );
  bc_pe bc_pe_884 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_884_clock),
    .reset(bc_pe_884_reset),
    .io_ho_input(bc_pe_884_io_ho_input),
    .io_ve_input(bc_pe_884_io_ve_input),
    .io_input_valid(bc_pe_884_io_input_valid),
    .io_iormac(bc_pe_884_io_iormac),
    .io_ve_out(bc_pe_884_io_ve_out),
    .io_ho_out(bc_pe_884_io_ho_out),
    .io_res_out(bc_pe_884_io_res_out)
  );
  bc_pe bc_pe_885 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_885_clock),
    .reset(bc_pe_885_reset),
    .io_ho_input(bc_pe_885_io_ho_input),
    .io_ve_input(bc_pe_885_io_ve_input),
    .io_input_valid(bc_pe_885_io_input_valid),
    .io_iormac(bc_pe_885_io_iormac),
    .io_ve_out(bc_pe_885_io_ve_out),
    .io_ho_out(bc_pe_885_io_ho_out),
    .io_res_out(bc_pe_885_io_res_out)
  );
  bc_pe bc_pe_886 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_886_clock),
    .reset(bc_pe_886_reset),
    .io_ho_input(bc_pe_886_io_ho_input),
    .io_ve_input(bc_pe_886_io_ve_input),
    .io_input_valid(bc_pe_886_io_input_valid),
    .io_iormac(bc_pe_886_io_iormac),
    .io_ve_out(bc_pe_886_io_ve_out),
    .io_ho_out(bc_pe_886_io_ho_out),
    .io_res_out(bc_pe_886_io_res_out)
  );
  bc_pe bc_pe_887 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_887_clock),
    .reset(bc_pe_887_reset),
    .io_ho_input(bc_pe_887_io_ho_input),
    .io_ve_input(bc_pe_887_io_ve_input),
    .io_input_valid(bc_pe_887_io_input_valid),
    .io_iormac(bc_pe_887_io_iormac),
    .io_ve_out(bc_pe_887_io_ve_out),
    .io_ho_out(bc_pe_887_io_ho_out),
    .io_res_out(bc_pe_887_io_res_out)
  );
  bc_pe bc_pe_888 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_888_clock),
    .reset(bc_pe_888_reset),
    .io_ho_input(bc_pe_888_io_ho_input),
    .io_ve_input(bc_pe_888_io_ve_input),
    .io_input_valid(bc_pe_888_io_input_valid),
    .io_iormac(bc_pe_888_io_iormac),
    .io_ve_out(bc_pe_888_io_ve_out),
    .io_ho_out(bc_pe_888_io_ho_out),
    .io_res_out(bc_pe_888_io_res_out)
  );
  bc_pe bc_pe_889 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_889_clock),
    .reset(bc_pe_889_reset),
    .io_ho_input(bc_pe_889_io_ho_input),
    .io_ve_input(bc_pe_889_io_ve_input),
    .io_input_valid(bc_pe_889_io_input_valid),
    .io_iormac(bc_pe_889_io_iormac),
    .io_ve_out(bc_pe_889_io_ve_out),
    .io_ho_out(bc_pe_889_io_ho_out),
    .io_res_out(bc_pe_889_io_res_out)
  );
  bc_pe bc_pe_890 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_890_clock),
    .reset(bc_pe_890_reset),
    .io_ho_input(bc_pe_890_io_ho_input),
    .io_ve_input(bc_pe_890_io_ve_input),
    .io_input_valid(bc_pe_890_io_input_valid),
    .io_iormac(bc_pe_890_io_iormac),
    .io_ve_out(bc_pe_890_io_ve_out),
    .io_ho_out(bc_pe_890_io_ho_out),
    .io_res_out(bc_pe_890_io_res_out)
  );
  bc_pe bc_pe_891 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_891_clock),
    .reset(bc_pe_891_reset),
    .io_ho_input(bc_pe_891_io_ho_input),
    .io_ve_input(bc_pe_891_io_ve_input),
    .io_input_valid(bc_pe_891_io_input_valid),
    .io_iormac(bc_pe_891_io_iormac),
    .io_ve_out(bc_pe_891_io_ve_out),
    .io_ho_out(bc_pe_891_io_ho_out),
    .io_res_out(bc_pe_891_io_res_out)
  );
  bc_pe bc_pe_892 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_892_clock),
    .reset(bc_pe_892_reset),
    .io_ho_input(bc_pe_892_io_ho_input),
    .io_ve_input(bc_pe_892_io_ve_input),
    .io_input_valid(bc_pe_892_io_input_valid),
    .io_iormac(bc_pe_892_io_iormac),
    .io_ve_out(bc_pe_892_io_ve_out),
    .io_ho_out(bc_pe_892_io_ho_out),
    .io_res_out(bc_pe_892_io_res_out)
  );
  bc_pe bc_pe_893 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_893_clock),
    .reset(bc_pe_893_reset),
    .io_ho_input(bc_pe_893_io_ho_input),
    .io_ve_input(bc_pe_893_io_ve_input),
    .io_input_valid(bc_pe_893_io_input_valid),
    .io_iormac(bc_pe_893_io_iormac),
    .io_ve_out(bc_pe_893_io_ve_out),
    .io_ho_out(bc_pe_893_io_ho_out),
    .io_res_out(bc_pe_893_io_res_out)
  );
  bc_pe bc_pe_894 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_894_clock),
    .reset(bc_pe_894_reset),
    .io_ho_input(bc_pe_894_io_ho_input),
    .io_ve_input(bc_pe_894_io_ve_input),
    .io_input_valid(bc_pe_894_io_input_valid),
    .io_iormac(bc_pe_894_io_iormac),
    .io_ve_out(bc_pe_894_io_ve_out),
    .io_ho_out(bc_pe_894_io_ho_out),
    .io_res_out(bc_pe_894_io_res_out)
  );
  bc_pe bc_pe_895 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_895_clock),
    .reset(bc_pe_895_reset),
    .io_ho_input(bc_pe_895_io_ho_input),
    .io_ve_input(bc_pe_895_io_ve_input),
    .io_input_valid(bc_pe_895_io_input_valid),
    .io_iormac(bc_pe_895_io_iormac),
    .io_ve_out(bc_pe_895_io_ve_out),
    .io_ho_out(bc_pe_895_io_ho_out),
    .io_res_out(bc_pe_895_io_res_out)
  );
  bc_pe bc_pe_896 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_896_clock),
    .reset(bc_pe_896_reset),
    .io_ho_input(bc_pe_896_io_ho_input),
    .io_ve_input(bc_pe_896_io_ve_input),
    .io_input_valid(bc_pe_896_io_input_valid),
    .io_iormac(bc_pe_896_io_iormac),
    .io_ve_out(bc_pe_896_io_ve_out),
    .io_ho_out(bc_pe_896_io_ho_out),
    .io_res_out(bc_pe_896_io_res_out)
  );
  bc_pe bc_pe_897 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_897_clock),
    .reset(bc_pe_897_reset),
    .io_ho_input(bc_pe_897_io_ho_input),
    .io_ve_input(bc_pe_897_io_ve_input),
    .io_input_valid(bc_pe_897_io_input_valid),
    .io_iormac(bc_pe_897_io_iormac),
    .io_ve_out(bc_pe_897_io_ve_out),
    .io_ho_out(bc_pe_897_io_ho_out),
    .io_res_out(bc_pe_897_io_res_out)
  );
  bc_pe bc_pe_898 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_898_clock),
    .reset(bc_pe_898_reset),
    .io_ho_input(bc_pe_898_io_ho_input),
    .io_ve_input(bc_pe_898_io_ve_input),
    .io_input_valid(bc_pe_898_io_input_valid),
    .io_iormac(bc_pe_898_io_iormac),
    .io_ve_out(bc_pe_898_io_ve_out),
    .io_ho_out(bc_pe_898_io_ho_out),
    .io_res_out(bc_pe_898_io_res_out)
  );
  bc_pe bc_pe_899 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_899_clock),
    .reset(bc_pe_899_reset),
    .io_ho_input(bc_pe_899_io_ho_input),
    .io_ve_input(bc_pe_899_io_ve_input),
    .io_input_valid(bc_pe_899_io_input_valid),
    .io_iormac(bc_pe_899_io_iormac),
    .io_ve_out(bc_pe_899_io_ve_out),
    .io_ho_out(bc_pe_899_io_ho_out),
    .io_res_out(bc_pe_899_io_res_out)
  );
  bc_pe bc_pe_900 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_900_clock),
    .reset(bc_pe_900_reset),
    .io_ho_input(bc_pe_900_io_ho_input),
    .io_ve_input(bc_pe_900_io_ve_input),
    .io_input_valid(bc_pe_900_io_input_valid),
    .io_iormac(bc_pe_900_io_iormac),
    .io_ve_out(bc_pe_900_io_ve_out),
    .io_ho_out(bc_pe_900_io_ho_out),
    .io_res_out(bc_pe_900_io_res_out)
  );
  bc_pe bc_pe_901 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_901_clock),
    .reset(bc_pe_901_reset),
    .io_ho_input(bc_pe_901_io_ho_input),
    .io_ve_input(bc_pe_901_io_ve_input),
    .io_input_valid(bc_pe_901_io_input_valid),
    .io_iormac(bc_pe_901_io_iormac),
    .io_ve_out(bc_pe_901_io_ve_out),
    .io_ho_out(bc_pe_901_io_ho_out),
    .io_res_out(bc_pe_901_io_res_out)
  );
  bc_pe bc_pe_902 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_902_clock),
    .reset(bc_pe_902_reset),
    .io_ho_input(bc_pe_902_io_ho_input),
    .io_ve_input(bc_pe_902_io_ve_input),
    .io_input_valid(bc_pe_902_io_input_valid),
    .io_iormac(bc_pe_902_io_iormac),
    .io_ve_out(bc_pe_902_io_ve_out),
    .io_ho_out(bc_pe_902_io_ho_out),
    .io_res_out(bc_pe_902_io_res_out)
  );
  bc_pe bc_pe_903 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_903_clock),
    .reset(bc_pe_903_reset),
    .io_ho_input(bc_pe_903_io_ho_input),
    .io_ve_input(bc_pe_903_io_ve_input),
    .io_input_valid(bc_pe_903_io_input_valid),
    .io_iormac(bc_pe_903_io_iormac),
    .io_ve_out(bc_pe_903_io_ve_out),
    .io_ho_out(bc_pe_903_io_ho_out),
    .io_res_out(bc_pe_903_io_res_out)
  );
  bc_pe bc_pe_904 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_904_clock),
    .reset(bc_pe_904_reset),
    .io_ho_input(bc_pe_904_io_ho_input),
    .io_ve_input(bc_pe_904_io_ve_input),
    .io_input_valid(bc_pe_904_io_input_valid),
    .io_iormac(bc_pe_904_io_iormac),
    .io_ve_out(bc_pe_904_io_ve_out),
    .io_ho_out(bc_pe_904_io_ho_out),
    .io_res_out(bc_pe_904_io_res_out)
  );
  bc_pe bc_pe_905 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_905_clock),
    .reset(bc_pe_905_reset),
    .io_ho_input(bc_pe_905_io_ho_input),
    .io_ve_input(bc_pe_905_io_ve_input),
    .io_input_valid(bc_pe_905_io_input_valid),
    .io_iormac(bc_pe_905_io_iormac),
    .io_ve_out(bc_pe_905_io_ve_out),
    .io_ho_out(bc_pe_905_io_ho_out),
    .io_res_out(bc_pe_905_io_res_out)
  );
  bc_pe bc_pe_906 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_906_clock),
    .reset(bc_pe_906_reset),
    .io_ho_input(bc_pe_906_io_ho_input),
    .io_ve_input(bc_pe_906_io_ve_input),
    .io_input_valid(bc_pe_906_io_input_valid),
    .io_iormac(bc_pe_906_io_iormac),
    .io_ve_out(bc_pe_906_io_ve_out),
    .io_ho_out(bc_pe_906_io_ho_out),
    .io_res_out(bc_pe_906_io_res_out)
  );
  bc_pe bc_pe_907 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_907_clock),
    .reset(bc_pe_907_reset),
    .io_ho_input(bc_pe_907_io_ho_input),
    .io_ve_input(bc_pe_907_io_ve_input),
    .io_input_valid(bc_pe_907_io_input_valid),
    .io_iormac(bc_pe_907_io_iormac),
    .io_ve_out(bc_pe_907_io_ve_out),
    .io_ho_out(bc_pe_907_io_ho_out),
    .io_res_out(bc_pe_907_io_res_out)
  );
  bc_pe bc_pe_908 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_908_clock),
    .reset(bc_pe_908_reset),
    .io_ho_input(bc_pe_908_io_ho_input),
    .io_ve_input(bc_pe_908_io_ve_input),
    .io_input_valid(bc_pe_908_io_input_valid),
    .io_iormac(bc_pe_908_io_iormac),
    .io_ve_out(bc_pe_908_io_ve_out),
    .io_ho_out(bc_pe_908_io_ho_out),
    .io_res_out(bc_pe_908_io_res_out)
  );
  bc_pe bc_pe_909 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_909_clock),
    .reset(bc_pe_909_reset),
    .io_ho_input(bc_pe_909_io_ho_input),
    .io_ve_input(bc_pe_909_io_ve_input),
    .io_input_valid(bc_pe_909_io_input_valid),
    .io_iormac(bc_pe_909_io_iormac),
    .io_ve_out(bc_pe_909_io_ve_out),
    .io_ho_out(bc_pe_909_io_ho_out),
    .io_res_out(bc_pe_909_io_res_out)
  );
  bc_pe bc_pe_910 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_910_clock),
    .reset(bc_pe_910_reset),
    .io_ho_input(bc_pe_910_io_ho_input),
    .io_ve_input(bc_pe_910_io_ve_input),
    .io_input_valid(bc_pe_910_io_input_valid),
    .io_iormac(bc_pe_910_io_iormac),
    .io_ve_out(bc_pe_910_io_ve_out),
    .io_ho_out(bc_pe_910_io_ho_out),
    .io_res_out(bc_pe_910_io_res_out)
  );
  bc_pe bc_pe_911 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_911_clock),
    .reset(bc_pe_911_reset),
    .io_ho_input(bc_pe_911_io_ho_input),
    .io_ve_input(bc_pe_911_io_ve_input),
    .io_input_valid(bc_pe_911_io_input_valid),
    .io_iormac(bc_pe_911_io_iormac),
    .io_ve_out(bc_pe_911_io_ve_out),
    .io_ho_out(bc_pe_911_io_ho_out),
    .io_res_out(bc_pe_911_io_res_out)
  );
  bc_pe bc_pe_912 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_912_clock),
    .reset(bc_pe_912_reset),
    .io_ho_input(bc_pe_912_io_ho_input),
    .io_ve_input(bc_pe_912_io_ve_input),
    .io_input_valid(bc_pe_912_io_input_valid),
    .io_iormac(bc_pe_912_io_iormac),
    .io_ve_out(bc_pe_912_io_ve_out),
    .io_ho_out(bc_pe_912_io_ho_out),
    .io_res_out(bc_pe_912_io_res_out)
  );
  bc_pe bc_pe_913 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_913_clock),
    .reset(bc_pe_913_reset),
    .io_ho_input(bc_pe_913_io_ho_input),
    .io_ve_input(bc_pe_913_io_ve_input),
    .io_input_valid(bc_pe_913_io_input_valid),
    .io_iormac(bc_pe_913_io_iormac),
    .io_ve_out(bc_pe_913_io_ve_out),
    .io_ho_out(bc_pe_913_io_ho_out),
    .io_res_out(bc_pe_913_io_res_out)
  );
  bc_pe bc_pe_914 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_914_clock),
    .reset(bc_pe_914_reset),
    .io_ho_input(bc_pe_914_io_ho_input),
    .io_ve_input(bc_pe_914_io_ve_input),
    .io_input_valid(bc_pe_914_io_input_valid),
    .io_iormac(bc_pe_914_io_iormac),
    .io_ve_out(bc_pe_914_io_ve_out),
    .io_ho_out(bc_pe_914_io_ho_out),
    .io_res_out(bc_pe_914_io_res_out)
  );
  bc_pe bc_pe_915 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_915_clock),
    .reset(bc_pe_915_reset),
    .io_ho_input(bc_pe_915_io_ho_input),
    .io_ve_input(bc_pe_915_io_ve_input),
    .io_input_valid(bc_pe_915_io_input_valid),
    .io_iormac(bc_pe_915_io_iormac),
    .io_ve_out(bc_pe_915_io_ve_out),
    .io_ho_out(bc_pe_915_io_ho_out),
    .io_res_out(bc_pe_915_io_res_out)
  );
  bc_pe bc_pe_916 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_916_clock),
    .reset(bc_pe_916_reset),
    .io_ho_input(bc_pe_916_io_ho_input),
    .io_ve_input(bc_pe_916_io_ve_input),
    .io_input_valid(bc_pe_916_io_input_valid),
    .io_iormac(bc_pe_916_io_iormac),
    .io_ve_out(bc_pe_916_io_ve_out),
    .io_ho_out(bc_pe_916_io_ho_out),
    .io_res_out(bc_pe_916_io_res_out)
  );
  bc_pe bc_pe_917 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_917_clock),
    .reset(bc_pe_917_reset),
    .io_ho_input(bc_pe_917_io_ho_input),
    .io_ve_input(bc_pe_917_io_ve_input),
    .io_input_valid(bc_pe_917_io_input_valid),
    .io_iormac(bc_pe_917_io_iormac),
    .io_ve_out(bc_pe_917_io_ve_out),
    .io_ho_out(bc_pe_917_io_ho_out),
    .io_res_out(bc_pe_917_io_res_out)
  );
  bc_pe bc_pe_918 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_918_clock),
    .reset(bc_pe_918_reset),
    .io_ho_input(bc_pe_918_io_ho_input),
    .io_ve_input(bc_pe_918_io_ve_input),
    .io_input_valid(bc_pe_918_io_input_valid),
    .io_iormac(bc_pe_918_io_iormac),
    .io_ve_out(bc_pe_918_io_ve_out),
    .io_ho_out(bc_pe_918_io_ho_out),
    .io_res_out(bc_pe_918_io_res_out)
  );
  bc_pe bc_pe_919 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_919_clock),
    .reset(bc_pe_919_reset),
    .io_ho_input(bc_pe_919_io_ho_input),
    .io_ve_input(bc_pe_919_io_ve_input),
    .io_input_valid(bc_pe_919_io_input_valid),
    .io_iormac(bc_pe_919_io_iormac),
    .io_ve_out(bc_pe_919_io_ve_out),
    .io_ho_out(bc_pe_919_io_ho_out),
    .io_res_out(bc_pe_919_io_res_out)
  );
  bc_pe bc_pe_920 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_920_clock),
    .reset(bc_pe_920_reset),
    .io_ho_input(bc_pe_920_io_ho_input),
    .io_ve_input(bc_pe_920_io_ve_input),
    .io_input_valid(bc_pe_920_io_input_valid),
    .io_iormac(bc_pe_920_io_iormac),
    .io_ve_out(bc_pe_920_io_ve_out),
    .io_ho_out(bc_pe_920_io_ho_out),
    .io_res_out(bc_pe_920_io_res_out)
  );
  bc_pe bc_pe_921 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_921_clock),
    .reset(bc_pe_921_reset),
    .io_ho_input(bc_pe_921_io_ho_input),
    .io_ve_input(bc_pe_921_io_ve_input),
    .io_input_valid(bc_pe_921_io_input_valid),
    .io_iormac(bc_pe_921_io_iormac),
    .io_ve_out(bc_pe_921_io_ve_out),
    .io_ho_out(bc_pe_921_io_ho_out),
    .io_res_out(bc_pe_921_io_res_out)
  );
  bc_pe bc_pe_922 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_922_clock),
    .reset(bc_pe_922_reset),
    .io_ho_input(bc_pe_922_io_ho_input),
    .io_ve_input(bc_pe_922_io_ve_input),
    .io_input_valid(bc_pe_922_io_input_valid),
    .io_iormac(bc_pe_922_io_iormac),
    .io_ve_out(bc_pe_922_io_ve_out),
    .io_ho_out(bc_pe_922_io_ho_out),
    .io_res_out(bc_pe_922_io_res_out)
  );
  bc_pe bc_pe_923 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_923_clock),
    .reset(bc_pe_923_reset),
    .io_ho_input(bc_pe_923_io_ho_input),
    .io_ve_input(bc_pe_923_io_ve_input),
    .io_input_valid(bc_pe_923_io_input_valid),
    .io_iormac(bc_pe_923_io_iormac),
    .io_ve_out(bc_pe_923_io_ve_out),
    .io_ho_out(bc_pe_923_io_ho_out),
    .io_res_out(bc_pe_923_io_res_out)
  );
  bc_pe bc_pe_924 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_924_clock),
    .reset(bc_pe_924_reset),
    .io_ho_input(bc_pe_924_io_ho_input),
    .io_ve_input(bc_pe_924_io_ve_input),
    .io_input_valid(bc_pe_924_io_input_valid),
    .io_iormac(bc_pe_924_io_iormac),
    .io_ve_out(bc_pe_924_io_ve_out),
    .io_ho_out(bc_pe_924_io_ho_out),
    .io_res_out(bc_pe_924_io_res_out)
  );
  bc_pe bc_pe_925 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_925_clock),
    .reset(bc_pe_925_reset),
    .io_ho_input(bc_pe_925_io_ho_input),
    .io_ve_input(bc_pe_925_io_ve_input),
    .io_input_valid(bc_pe_925_io_input_valid),
    .io_iormac(bc_pe_925_io_iormac),
    .io_ve_out(bc_pe_925_io_ve_out),
    .io_ho_out(bc_pe_925_io_ho_out),
    .io_res_out(bc_pe_925_io_res_out)
  );
  bc_pe bc_pe_926 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_926_clock),
    .reset(bc_pe_926_reset),
    .io_ho_input(bc_pe_926_io_ho_input),
    .io_ve_input(bc_pe_926_io_ve_input),
    .io_input_valid(bc_pe_926_io_input_valid),
    .io_iormac(bc_pe_926_io_iormac),
    .io_ve_out(bc_pe_926_io_ve_out),
    .io_ho_out(bc_pe_926_io_ho_out),
    .io_res_out(bc_pe_926_io_res_out)
  );
  bc_pe bc_pe_927 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_927_clock),
    .reset(bc_pe_927_reset),
    .io_ho_input(bc_pe_927_io_ho_input),
    .io_ve_input(bc_pe_927_io_ve_input),
    .io_input_valid(bc_pe_927_io_input_valid),
    .io_iormac(bc_pe_927_io_iormac),
    .io_ve_out(bc_pe_927_io_ve_out),
    .io_ho_out(bc_pe_927_io_ho_out),
    .io_res_out(bc_pe_927_io_res_out)
  );
  bc_pe bc_pe_928 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_928_clock),
    .reset(bc_pe_928_reset),
    .io_ho_input(bc_pe_928_io_ho_input),
    .io_ve_input(bc_pe_928_io_ve_input),
    .io_input_valid(bc_pe_928_io_input_valid),
    .io_iormac(bc_pe_928_io_iormac),
    .io_ve_out(bc_pe_928_io_ve_out),
    .io_ho_out(bc_pe_928_io_ho_out),
    .io_res_out(bc_pe_928_io_res_out)
  );
  bc_pe bc_pe_929 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_929_clock),
    .reset(bc_pe_929_reset),
    .io_ho_input(bc_pe_929_io_ho_input),
    .io_ve_input(bc_pe_929_io_ve_input),
    .io_input_valid(bc_pe_929_io_input_valid),
    .io_iormac(bc_pe_929_io_iormac),
    .io_ve_out(bc_pe_929_io_ve_out),
    .io_ho_out(bc_pe_929_io_ho_out),
    .io_res_out(bc_pe_929_io_res_out)
  );
  bc_pe bc_pe_930 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_930_clock),
    .reset(bc_pe_930_reset),
    .io_ho_input(bc_pe_930_io_ho_input),
    .io_ve_input(bc_pe_930_io_ve_input),
    .io_input_valid(bc_pe_930_io_input_valid),
    .io_iormac(bc_pe_930_io_iormac),
    .io_ve_out(bc_pe_930_io_ve_out),
    .io_ho_out(bc_pe_930_io_ho_out),
    .io_res_out(bc_pe_930_io_res_out)
  );
  bc_pe bc_pe_931 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_931_clock),
    .reset(bc_pe_931_reset),
    .io_ho_input(bc_pe_931_io_ho_input),
    .io_ve_input(bc_pe_931_io_ve_input),
    .io_input_valid(bc_pe_931_io_input_valid),
    .io_iormac(bc_pe_931_io_iormac),
    .io_ve_out(bc_pe_931_io_ve_out),
    .io_ho_out(bc_pe_931_io_ho_out),
    .io_res_out(bc_pe_931_io_res_out)
  );
  bc_pe bc_pe_932 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_932_clock),
    .reset(bc_pe_932_reset),
    .io_ho_input(bc_pe_932_io_ho_input),
    .io_ve_input(bc_pe_932_io_ve_input),
    .io_input_valid(bc_pe_932_io_input_valid),
    .io_iormac(bc_pe_932_io_iormac),
    .io_ve_out(bc_pe_932_io_ve_out),
    .io_ho_out(bc_pe_932_io_ho_out),
    .io_res_out(bc_pe_932_io_res_out)
  );
  bc_pe bc_pe_933 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_933_clock),
    .reset(bc_pe_933_reset),
    .io_ho_input(bc_pe_933_io_ho_input),
    .io_ve_input(bc_pe_933_io_ve_input),
    .io_input_valid(bc_pe_933_io_input_valid),
    .io_iormac(bc_pe_933_io_iormac),
    .io_ve_out(bc_pe_933_io_ve_out),
    .io_ho_out(bc_pe_933_io_ho_out),
    .io_res_out(bc_pe_933_io_res_out)
  );
  bc_pe bc_pe_934 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_934_clock),
    .reset(bc_pe_934_reset),
    .io_ho_input(bc_pe_934_io_ho_input),
    .io_ve_input(bc_pe_934_io_ve_input),
    .io_input_valid(bc_pe_934_io_input_valid),
    .io_iormac(bc_pe_934_io_iormac),
    .io_ve_out(bc_pe_934_io_ve_out),
    .io_ho_out(bc_pe_934_io_ho_out),
    .io_res_out(bc_pe_934_io_res_out)
  );
  bc_pe bc_pe_935 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_935_clock),
    .reset(bc_pe_935_reset),
    .io_ho_input(bc_pe_935_io_ho_input),
    .io_ve_input(bc_pe_935_io_ve_input),
    .io_input_valid(bc_pe_935_io_input_valid),
    .io_iormac(bc_pe_935_io_iormac),
    .io_ve_out(bc_pe_935_io_ve_out),
    .io_ho_out(bc_pe_935_io_ho_out),
    .io_res_out(bc_pe_935_io_res_out)
  );
  bc_pe bc_pe_936 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_936_clock),
    .reset(bc_pe_936_reset),
    .io_ho_input(bc_pe_936_io_ho_input),
    .io_ve_input(bc_pe_936_io_ve_input),
    .io_input_valid(bc_pe_936_io_input_valid),
    .io_iormac(bc_pe_936_io_iormac),
    .io_ve_out(bc_pe_936_io_ve_out),
    .io_ho_out(bc_pe_936_io_ho_out),
    .io_res_out(bc_pe_936_io_res_out)
  );
  bc_pe bc_pe_937 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_937_clock),
    .reset(bc_pe_937_reset),
    .io_ho_input(bc_pe_937_io_ho_input),
    .io_ve_input(bc_pe_937_io_ve_input),
    .io_input_valid(bc_pe_937_io_input_valid),
    .io_iormac(bc_pe_937_io_iormac),
    .io_ve_out(bc_pe_937_io_ve_out),
    .io_ho_out(bc_pe_937_io_ho_out),
    .io_res_out(bc_pe_937_io_res_out)
  );
  bc_pe bc_pe_938 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_938_clock),
    .reset(bc_pe_938_reset),
    .io_ho_input(bc_pe_938_io_ho_input),
    .io_ve_input(bc_pe_938_io_ve_input),
    .io_input_valid(bc_pe_938_io_input_valid),
    .io_iormac(bc_pe_938_io_iormac),
    .io_ve_out(bc_pe_938_io_ve_out),
    .io_ho_out(bc_pe_938_io_ho_out),
    .io_res_out(bc_pe_938_io_res_out)
  );
  bc_pe bc_pe_939 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_939_clock),
    .reset(bc_pe_939_reset),
    .io_ho_input(bc_pe_939_io_ho_input),
    .io_ve_input(bc_pe_939_io_ve_input),
    .io_input_valid(bc_pe_939_io_input_valid),
    .io_iormac(bc_pe_939_io_iormac),
    .io_ve_out(bc_pe_939_io_ve_out),
    .io_ho_out(bc_pe_939_io_ho_out),
    .io_res_out(bc_pe_939_io_res_out)
  );
  bc_pe bc_pe_940 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_940_clock),
    .reset(bc_pe_940_reset),
    .io_ho_input(bc_pe_940_io_ho_input),
    .io_ve_input(bc_pe_940_io_ve_input),
    .io_input_valid(bc_pe_940_io_input_valid),
    .io_iormac(bc_pe_940_io_iormac),
    .io_ve_out(bc_pe_940_io_ve_out),
    .io_ho_out(bc_pe_940_io_ho_out),
    .io_res_out(bc_pe_940_io_res_out)
  );
  bc_pe bc_pe_941 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_941_clock),
    .reset(bc_pe_941_reset),
    .io_ho_input(bc_pe_941_io_ho_input),
    .io_ve_input(bc_pe_941_io_ve_input),
    .io_input_valid(bc_pe_941_io_input_valid),
    .io_iormac(bc_pe_941_io_iormac),
    .io_ve_out(bc_pe_941_io_ve_out),
    .io_ho_out(bc_pe_941_io_ho_out),
    .io_res_out(bc_pe_941_io_res_out)
  );
  bc_pe bc_pe_942 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_942_clock),
    .reset(bc_pe_942_reset),
    .io_ho_input(bc_pe_942_io_ho_input),
    .io_ve_input(bc_pe_942_io_ve_input),
    .io_input_valid(bc_pe_942_io_input_valid),
    .io_iormac(bc_pe_942_io_iormac),
    .io_ve_out(bc_pe_942_io_ve_out),
    .io_ho_out(bc_pe_942_io_ho_out),
    .io_res_out(bc_pe_942_io_res_out)
  );
  bc_pe bc_pe_943 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_943_clock),
    .reset(bc_pe_943_reset),
    .io_ho_input(bc_pe_943_io_ho_input),
    .io_ve_input(bc_pe_943_io_ve_input),
    .io_input_valid(bc_pe_943_io_input_valid),
    .io_iormac(bc_pe_943_io_iormac),
    .io_ve_out(bc_pe_943_io_ve_out),
    .io_ho_out(bc_pe_943_io_ho_out),
    .io_res_out(bc_pe_943_io_res_out)
  );
  bc_pe bc_pe_944 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_944_clock),
    .reset(bc_pe_944_reset),
    .io_ho_input(bc_pe_944_io_ho_input),
    .io_ve_input(bc_pe_944_io_ve_input),
    .io_input_valid(bc_pe_944_io_input_valid),
    .io_iormac(bc_pe_944_io_iormac),
    .io_ve_out(bc_pe_944_io_ve_out),
    .io_ho_out(bc_pe_944_io_ho_out),
    .io_res_out(bc_pe_944_io_res_out)
  );
  bc_pe bc_pe_945 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_945_clock),
    .reset(bc_pe_945_reset),
    .io_ho_input(bc_pe_945_io_ho_input),
    .io_ve_input(bc_pe_945_io_ve_input),
    .io_input_valid(bc_pe_945_io_input_valid),
    .io_iormac(bc_pe_945_io_iormac),
    .io_ve_out(bc_pe_945_io_ve_out),
    .io_ho_out(bc_pe_945_io_ho_out),
    .io_res_out(bc_pe_945_io_res_out)
  );
  bc_pe bc_pe_946 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_946_clock),
    .reset(bc_pe_946_reset),
    .io_ho_input(bc_pe_946_io_ho_input),
    .io_ve_input(bc_pe_946_io_ve_input),
    .io_input_valid(bc_pe_946_io_input_valid),
    .io_iormac(bc_pe_946_io_iormac),
    .io_ve_out(bc_pe_946_io_ve_out),
    .io_ho_out(bc_pe_946_io_ho_out),
    .io_res_out(bc_pe_946_io_res_out)
  );
  bc_pe bc_pe_947 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_947_clock),
    .reset(bc_pe_947_reset),
    .io_ho_input(bc_pe_947_io_ho_input),
    .io_ve_input(bc_pe_947_io_ve_input),
    .io_input_valid(bc_pe_947_io_input_valid),
    .io_iormac(bc_pe_947_io_iormac),
    .io_ve_out(bc_pe_947_io_ve_out),
    .io_ho_out(bc_pe_947_io_ho_out),
    .io_res_out(bc_pe_947_io_res_out)
  );
  bc_pe bc_pe_948 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_948_clock),
    .reset(bc_pe_948_reset),
    .io_ho_input(bc_pe_948_io_ho_input),
    .io_ve_input(bc_pe_948_io_ve_input),
    .io_input_valid(bc_pe_948_io_input_valid),
    .io_iormac(bc_pe_948_io_iormac),
    .io_ve_out(bc_pe_948_io_ve_out),
    .io_ho_out(bc_pe_948_io_ho_out),
    .io_res_out(bc_pe_948_io_res_out)
  );
  bc_pe bc_pe_949 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_949_clock),
    .reset(bc_pe_949_reset),
    .io_ho_input(bc_pe_949_io_ho_input),
    .io_ve_input(bc_pe_949_io_ve_input),
    .io_input_valid(bc_pe_949_io_input_valid),
    .io_iormac(bc_pe_949_io_iormac),
    .io_ve_out(bc_pe_949_io_ve_out),
    .io_ho_out(bc_pe_949_io_ho_out),
    .io_res_out(bc_pe_949_io_res_out)
  );
  bc_pe bc_pe_950 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_950_clock),
    .reset(bc_pe_950_reset),
    .io_ho_input(bc_pe_950_io_ho_input),
    .io_ve_input(bc_pe_950_io_ve_input),
    .io_input_valid(bc_pe_950_io_input_valid),
    .io_iormac(bc_pe_950_io_iormac),
    .io_ve_out(bc_pe_950_io_ve_out),
    .io_ho_out(bc_pe_950_io_ho_out),
    .io_res_out(bc_pe_950_io_res_out)
  );
  bc_pe bc_pe_951 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_951_clock),
    .reset(bc_pe_951_reset),
    .io_ho_input(bc_pe_951_io_ho_input),
    .io_ve_input(bc_pe_951_io_ve_input),
    .io_input_valid(bc_pe_951_io_input_valid),
    .io_iormac(bc_pe_951_io_iormac),
    .io_ve_out(bc_pe_951_io_ve_out),
    .io_ho_out(bc_pe_951_io_ho_out),
    .io_res_out(bc_pe_951_io_res_out)
  );
  bc_pe bc_pe_952 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_952_clock),
    .reset(bc_pe_952_reset),
    .io_ho_input(bc_pe_952_io_ho_input),
    .io_ve_input(bc_pe_952_io_ve_input),
    .io_input_valid(bc_pe_952_io_input_valid),
    .io_iormac(bc_pe_952_io_iormac),
    .io_ve_out(bc_pe_952_io_ve_out),
    .io_ho_out(bc_pe_952_io_ho_out),
    .io_res_out(bc_pe_952_io_res_out)
  );
  bc_pe bc_pe_953 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_953_clock),
    .reset(bc_pe_953_reset),
    .io_ho_input(bc_pe_953_io_ho_input),
    .io_ve_input(bc_pe_953_io_ve_input),
    .io_input_valid(bc_pe_953_io_input_valid),
    .io_iormac(bc_pe_953_io_iormac),
    .io_ve_out(bc_pe_953_io_ve_out),
    .io_ho_out(bc_pe_953_io_ho_out),
    .io_res_out(bc_pe_953_io_res_out)
  );
  bc_pe bc_pe_954 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_954_clock),
    .reset(bc_pe_954_reset),
    .io_ho_input(bc_pe_954_io_ho_input),
    .io_ve_input(bc_pe_954_io_ve_input),
    .io_input_valid(bc_pe_954_io_input_valid),
    .io_iormac(bc_pe_954_io_iormac),
    .io_ve_out(bc_pe_954_io_ve_out),
    .io_ho_out(bc_pe_954_io_ho_out),
    .io_res_out(bc_pe_954_io_res_out)
  );
  bc_pe bc_pe_955 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_955_clock),
    .reset(bc_pe_955_reset),
    .io_ho_input(bc_pe_955_io_ho_input),
    .io_ve_input(bc_pe_955_io_ve_input),
    .io_input_valid(bc_pe_955_io_input_valid),
    .io_iormac(bc_pe_955_io_iormac),
    .io_ve_out(bc_pe_955_io_ve_out),
    .io_ho_out(bc_pe_955_io_ho_out),
    .io_res_out(bc_pe_955_io_res_out)
  );
  bc_pe bc_pe_956 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_956_clock),
    .reset(bc_pe_956_reset),
    .io_ho_input(bc_pe_956_io_ho_input),
    .io_ve_input(bc_pe_956_io_ve_input),
    .io_input_valid(bc_pe_956_io_input_valid),
    .io_iormac(bc_pe_956_io_iormac),
    .io_ve_out(bc_pe_956_io_ve_out),
    .io_ho_out(bc_pe_956_io_ho_out),
    .io_res_out(bc_pe_956_io_res_out)
  );
  bc_pe bc_pe_957 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_957_clock),
    .reset(bc_pe_957_reset),
    .io_ho_input(bc_pe_957_io_ho_input),
    .io_ve_input(bc_pe_957_io_ve_input),
    .io_input_valid(bc_pe_957_io_input_valid),
    .io_iormac(bc_pe_957_io_iormac),
    .io_ve_out(bc_pe_957_io_ve_out),
    .io_ho_out(bc_pe_957_io_ho_out),
    .io_res_out(bc_pe_957_io_res_out)
  );
  bc_pe bc_pe_958 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_958_clock),
    .reset(bc_pe_958_reset),
    .io_ho_input(bc_pe_958_io_ho_input),
    .io_ve_input(bc_pe_958_io_ve_input),
    .io_input_valid(bc_pe_958_io_input_valid),
    .io_iormac(bc_pe_958_io_iormac),
    .io_ve_out(bc_pe_958_io_ve_out),
    .io_ho_out(bc_pe_958_io_ho_out),
    .io_res_out(bc_pe_958_io_res_out)
  );
  bc_pe bc_pe_959 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_959_clock),
    .reset(bc_pe_959_reset),
    .io_ho_input(bc_pe_959_io_ho_input),
    .io_ve_input(bc_pe_959_io_ve_input),
    .io_input_valid(bc_pe_959_io_input_valid),
    .io_iormac(bc_pe_959_io_iormac),
    .io_ve_out(bc_pe_959_io_ve_out),
    .io_ho_out(bc_pe_959_io_ho_out),
    .io_res_out(bc_pe_959_io_res_out)
  );
  bc_pe bc_pe_960 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_960_clock),
    .reset(bc_pe_960_reset),
    .io_ho_input(bc_pe_960_io_ho_input),
    .io_ve_input(bc_pe_960_io_ve_input),
    .io_input_valid(bc_pe_960_io_input_valid),
    .io_iormac(bc_pe_960_io_iormac),
    .io_ve_out(bc_pe_960_io_ve_out),
    .io_ho_out(bc_pe_960_io_ho_out),
    .io_res_out(bc_pe_960_io_res_out)
  );
  bc_pe bc_pe_961 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_961_clock),
    .reset(bc_pe_961_reset),
    .io_ho_input(bc_pe_961_io_ho_input),
    .io_ve_input(bc_pe_961_io_ve_input),
    .io_input_valid(bc_pe_961_io_input_valid),
    .io_iormac(bc_pe_961_io_iormac),
    .io_ve_out(bc_pe_961_io_ve_out),
    .io_ho_out(bc_pe_961_io_ho_out),
    .io_res_out(bc_pe_961_io_res_out)
  );
  bc_pe bc_pe_962 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_962_clock),
    .reset(bc_pe_962_reset),
    .io_ho_input(bc_pe_962_io_ho_input),
    .io_ve_input(bc_pe_962_io_ve_input),
    .io_input_valid(bc_pe_962_io_input_valid),
    .io_iormac(bc_pe_962_io_iormac),
    .io_ve_out(bc_pe_962_io_ve_out),
    .io_ho_out(bc_pe_962_io_ho_out),
    .io_res_out(bc_pe_962_io_res_out)
  );
  bc_pe bc_pe_963 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_963_clock),
    .reset(bc_pe_963_reset),
    .io_ho_input(bc_pe_963_io_ho_input),
    .io_ve_input(bc_pe_963_io_ve_input),
    .io_input_valid(bc_pe_963_io_input_valid),
    .io_iormac(bc_pe_963_io_iormac),
    .io_ve_out(bc_pe_963_io_ve_out),
    .io_ho_out(bc_pe_963_io_ho_out),
    .io_res_out(bc_pe_963_io_res_out)
  );
  bc_pe bc_pe_964 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_964_clock),
    .reset(bc_pe_964_reset),
    .io_ho_input(bc_pe_964_io_ho_input),
    .io_ve_input(bc_pe_964_io_ve_input),
    .io_input_valid(bc_pe_964_io_input_valid),
    .io_iormac(bc_pe_964_io_iormac),
    .io_ve_out(bc_pe_964_io_ve_out),
    .io_ho_out(bc_pe_964_io_ho_out),
    .io_res_out(bc_pe_964_io_res_out)
  );
  bc_pe bc_pe_965 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_965_clock),
    .reset(bc_pe_965_reset),
    .io_ho_input(bc_pe_965_io_ho_input),
    .io_ve_input(bc_pe_965_io_ve_input),
    .io_input_valid(bc_pe_965_io_input_valid),
    .io_iormac(bc_pe_965_io_iormac),
    .io_ve_out(bc_pe_965_io_ve_out),
    .io_ho_out(bc_pe_965_io_ho_out),
    .io_res_out(bc_pe_965_io_res_out)
  );
  bc_pe bc_pe_966 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_966_clock),
    .reset(bc_pe_966_reset),
    .io_ho_input(bc_pe_966_io_ho_input),
    .io_ve_input(bc_pe_966_io_ve_input),
    .io_input_valid(bc_pe_966_io_input_valid),
    .io_iormac(bc_pe_966_io_iormac),
    .io_ve_out(bc_pe_966_io_ve_out),
    .io_ho_out(bc_pe_966_io_ho_out),
    .io_res_out(bc_pe_966_io_res_out)
  );
  bc_pe bc_pe_967 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_967_clock),
    .reset(bc_pe_967_reset),
    .io_ho_input(bc_pe_967_io_ho_input),
    .io_ve_input(bc_pe_967_io_ve_input),
    .io_input_valid(bc_pe_967_io_input_valid),
    .io_iormac(bc_pe_967_io_iormac),
    .io_ve_out(bc_pe_967_io_ve_out),
    .io_ho_out(bc_pe_967_io_ho_out),
    .io_res_out(bc_pe_967_io_res_out)
  );
  bc_pe bc_pe_968 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_968_clock),
    .reset(bc_pe_968_reset),
    .io_ho_input(bc_pe_968_io_ho_input),
    .io_ve_input(bc_pe_968_io_ve_input),
    .io_input_valid(bc_pe_968_io_input_valid),
    .io_iormac(bc_pe_968_io_iormac),
    .io_ve_out(bc_pe_968_io_ve_out),
    .io_ho_out(bc_pe_968_io_ho_out),
    .io_res_out(bc_pe_968_io_res_out)
  );
  bc_pe bc_pe_969 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_969_clock),
    .reset(bc_pe_969_reset),
    .io_ho_input(bc_pe_969_io_ho_input),
    .io_ve_input(bc_pe_969_io_ve_input),
    .io_input_valid(bc_pe_969_io_input_valid),
    .io_iormac(bc_pe_969_io_iormac),
    .io_ve_out(bc_pe_969_io_ve_out),
    .io_ho_out(bc_pe_969_io_ho_out),
    .io_res_out(bc_pe_969_io_res_out)
  );
  bc_pe bc_pe_970 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_970_clock),
    .reset(bc_pe_970_reset),
    .io_ho_input(bc_pe_970_io_ho_input),
    .io_ve_input(bc_pe_970_io_ve_input),
    .io_input_valid(bc_pe_970_io_input_valid),
    .io_iormac(bc_pe_970_io_iormac),
    .io_ve_out(bc_pe_970_io_ve_out),
    .io_ho_out(bc_pe_970_io_ho_out),
    .io_res_out(bc_pe_970_io_res_out)
  );
  bc_pe bc_pe_971 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_971_clock),
    .reset(bc_pe_971_reset),
    .io_ho_input(bc_pe_971_io_ho_input),
    .io_ve_input(bc_pe_971_io_ve_input),
    .io_input_valid(bc_pe_971_io_input_valid),
    .io_iormac(bc_pe_971_io_iormac),
    .io_ve_out(bc_pe_971_io_ve_out),
    .io_ho_out(bc_pe_971_io_ho_out),
    .io_res_out(bc_pe_971_io_res_out)
  );
  bc_pe bc_pe_972 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_972_clock),
    .reset(bc_pe_972_reset),
    .io_ho_input(bc_pe_972_io_ho_input),
    .io_ve_input(bc_pe_972_io_ve_input),
    .io_input_valid(bc_pe_972_io_input_valid),
    .io_iormac(bc_pe_972_io_iormac),
    .io_ve_out(bc_pe_972_io_ve_out),
    .io_ho_out(bc_pe_972_io_ho_out),
    .io_res_out(bc_pe_972_io_res_out)
  );
  bc_pe bc_pe_973 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_973_clock),
    .reset(bc_pe_973_reset),
    .io_ho_input(bc_pe_973_io_ho_input),
    .io_ve_input(bc_pe_973_io_ve_input),
    .io_input_valid(bc_pe_973_io_input_valid),
    .io_iormac(bc_pe_973_io_iormac),
    .io_ve_out(bc_pe_973_io_ve_out),
    .io_ho_out(bc_pe_973_io_ho_out),
    .io_res_out(bc_pe_973_io_res_out)
  );
  bc_pe bc_pe_974 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_974_clock),
    .reset(bc_pe_974_reset),
    .io_ho_input(bc_pe_974_io_ho_input),
    .io_ve_input(bc_pe_974_io_ve_input),
    .io_input_valid(bc_pe_974_io_input_valid),
    .io_iormac(bc_pe_974_io_iormac),
    .io_ve_out(bc_pe_974_io_ve_out),
    .io_ho_out(bc_pe_974_io_ho_out),
    .io_res_out(bc_pe_974_io_res_out)
  );
  bc_pe bc_pe_975 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_975_clock),
    .reset(bc_pe_975_reset),
    .io_ho_input(bc_pe_975_io_ho_input),
    .io_ve_input(bc_pe_975_io_ve_input),
    .io_input_valid(bc_pe_975_io_input_valid),
    .io_iormac(bc_pe_975_io_iormac),
    .io_ve_out(bc_pe_975_io_ve_out),
    .io_ho_out(bc_pe_975_io_ho_out),
    .io_res_out(bc_pe_975_io_res_out)
  );
  bc_pe bc_pe_976 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_976_clock),
    .reset(bc_pe_976_reset),
    .io_ho_input(bc_pe_976_io_ho_input),
    .io_ve_input(bc_pe_976_io_ve_input),
    .io_input_valid(bc_pe_976_io_input_valid),
    .io_iormac(bc_pe_976_io_iormac),
    .io_ve_out(bc_pe_976_io_ve_out),
    .io_ho_out(bc_pe_976_io_ho_out),
    .io_res_out(bc_pe_976_io_res_out)
  );
  bc_pe bc_pe_977 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_977_clock),
    .reset(bc_pe_977_reset),
    .io_ho_input(bc_pe_977_io_ho_input),
    .io_ve_input(bc_pe_977_io_ve_input),
    .io_input_valid(bc_pe_977_io_input_valid),
    .io_iormac(bc_pe_977_io_iormac),
    .io_ve_out(bc_pe_977_io_ve_out),
    .io_ho_out(bc_pe_977_io_ho_out),
    .io_res_out(bc_pe_977_io_res_out)
  );
  bc_pe bc_pe_978 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_978_clock),
    .reset(bc_pe_978_reset),
    .io_ho_input(bc_pe_978_io_ho_input),
    .io_ve_input(bc_pe_978_io_ve_input),
    .io_input_valid(bc_pe_978_io_input_valid),
    .io_iormac(bc_pe_978_io_iormac),
    .io_ve_out(bc_pe_978_io_ve_out),
    .io_ho_out(bc_pe_978_io_ho_out),
    .io_res_out(bc_pe_978_io_res_out)
  );
  bc_pe bc_pe_979 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_979_clock),
    .reset(bc_pe_979_reset),
    .io_ho_input(bc_pe_979_io_ho_input),
    .io_ve_input(bc_pe_979_io_ve_input),
    .io_input_valid(bc_pe_979_io_input_valid),
    .io_iormac(bc_pe_979_io_iormac),
    .io_ve_out(bc_pe_979_io_ve_out),
    .io_ho_out(bc_pe_979_io_ho_out),
    .io_res_out(bc_pe_979_io_res_out)
  );
  bc_pe bc_pe_980 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_980_clock),
    .reset(bc_pe_980_reset),
    .io_ho_input(bc_pe_980_io_ho_input),
    .io_ve_input(bc_pe_980_io_ve_input),
    .io_input_valid(bc_pe_980_io_input_valid),
    .io_iormac(bc_pe_980_io_iormac),
    .io_ve_out(bc_pe_980_io_ve_out),
    .io_ho_out(bc_pe_980_io_ho_out),
    .io_res_out(bc_pe_980_io_res_out)
  );
  bc_pe bc_pe_981 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_981_clock),
    .reset(bc_pe_981_reset),
    .io_ho_input(bc_pe_981_io_ho_input),
    .io_ve_input(bc_pe_981_io_ve_input),
    .io_input_valid(bc_pe_981_io_input_valid),
    .io_iormac(bc_pe_981_io_iormac),
    .io_ve_out(bc_pe_981_io_ve_out),
    .io_ho_out(bc_pe_981_io_ho_out),
    .io_res_out(bc_pe_981_io_res_out)
  );
  bc_pe bc_pe_982 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_982_clock),
    .reset(bc_pe_982_reset),
    .io_ho_input(bc_pe_982_io_ho_input),
    .io_ve_input(bc_pe_982_io_ve_input),
    .io_input_valid(bc_pe_982_io_input_valid),
    .io_iormac(bc_pe_982_io_iormac),
    .io_ve_out(bc_pe_982_io_ve_out),
    .io_ho_out(bc_pe_982_io_ho_out),
    .io_res_out(bc_pe_982_io_res_out)
  );
  bc_pe bc_pe_983 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_983_clock),
    .reset(bc_pe_983_reset),
    .io_ho_input(bc_pe_983_io_ho_input),
    .io_ve_input(bc_pe_983_io_ve_input),
    .io_input_valid(bc_pe_983_io_input_valid),
    .io_iormac(bc_pe_983_io_iormac),
    .io_ve_out(bc_pe_983_io_ve_out),
    .io_ho_out(bc_pe_983_io_ho_out),
    .io_res_out(bc_pe_983_io_res_out)
  );
  bc_pe bc_pe_984 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_984_clock),
    .reset(bc_pe_984_reset),
    .io_ho_input(bc_pe_984_io_ho_input),
    .io_ve_input(bc_pe_984_io_ve_input),
    .io_input_valid(bc_pe_984_io_input_valid),
    .io_iormac(bc_pe_984_io_iormac),
    .io_ve_out(bc_pe_984_io_ve_out),
    .io_ho_out(bc_pe_984_io_ho_out),
    .io_res_out(bc_pe_984_io_res_out)
  );
  bc_pe bc_pe_985 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_985_clock),
    .reset(bc_pe_985_reset),
    .io_ho_input(bc_pe_985_io_ho_input),
    .io_ve_input(bc_pe_985_io_ve_input),
    .io_input_valid(bc_pe_985_io_input_valid),
    .io_iormac(bc_pe_985_io_iormac),
    .io_ve_out(bc_pe_985_io_ve_out),
    .io_ho_out(bc_pe_985_io_ho_out),
    .io_res_out(bc_pe_985_io_res_out)
  );
  bc_pe bc_pe_986 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_986_clock),
    .reset(bc_pe_986_reset),
    .io_ho_input(bc_pe_986_io_ho_input),
    .io_ve_input(bc_pe_986_io_ve_input),
    .io_input_valid(bc_pe_986_io_input_valid),
    .io_iormac(bc_pe_986_io_iormac),
    .io_ve_out(bc_pe_986_io_ve_out),
    .io_ho_out(bc_pe_986_io_ho_out),
    .io_res_out(bc_pe_986_io_res_out)
  );
  bc_pe bc_pe_987 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_987_clock),
    .reset(bc_pe_987_reset),
    .io_ho_input(bc_pe_987_io_ho_input),
    .io_ve_input(bc_pe_987_io_ve_input),
    .io_input_valid(bc_pe_987_io_input_valid),
    .io_iormac(bc_pe_987_io_iormac),
    .io_ve_out(bc_pe_987_io_ve_out),
    .io_ho_out(bc_pe_987_io_ho_out),
    .io_res_out(bc_pe_987_io_res_out)
  );
  bc_pe bc_pe_988 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_988_clock),
    .reset(bc_pe_988_reset),
    .io_ho_input(bc_pe_988_io_ho_input),
    .io_ve_input(bc_pe_988_io_ve_input),
    .io_input_valid(bc_pe_988_io_input_valid),
    .io_iormac(bc_pe_988_io_iormac),
    .io_ve_out(bc_pe_988_io_ve_out),
    .io_ho_out(bc_pe_988_io_ho_out),
    .io_res_out(bc_pe_988_io_res_out)
  );
  bc_pe bc_pe_989 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_989_clock),
    .reset(bc_pe_989_reset),
    .io_ho_input(bc_pe_989_io_ho_input),
    .io_ve_input(bc_pe_989_io_ve_input),
    .io_input_valid(bc_pe_989_io_input_valid),
    .io_iormac(bc_pe_989_io_iormac),
    .io_ve_out(bc_pe_989_io_ve_out),
    .io_ho_out(bc_pe_989_io_ho_out),
    .io_res_out(bc_pe_989_io_res_out)
  );
  bc_pe bc_pe_990 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_990_clock),
    .reset(bc_pe_990_reset),
    .io_ho_input(bc_pe_990_io_ho_input),
    .io_ve_input(bc_pe_990_io_ve_input),
    .io_input_valid(bc_pe_990_io_input_valid),
    .io_iormac(bc_pe_990_io_iormac),
    .io_ve_out(bc_pe_990_io_ve_out),
    .io_ho_out(bc_pe_990_io_ho_out),
    .io_res_out(bc_pe_990_io_res_out)
  );
  bc_pe bc_pe_991 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_991_clock),
    .reset(bc_pe_991_reset),
    .io_ho_input(bc_pe_991_io_ho_input),
    .io_ve_input(bc_pe_991_io_ve_input),
    .io_input_valid(bc_pe_991_io_input_valid),
    .io_iormac(bc_pe_991_io_iormac),
    .io_ve_out(bc_pe_991_io_ve_out),
    .io_ho_out(bc_pe_991_io_ho_out),
    .io_res_out(bc_pe_991_io_res_out)
  );
  bc_pe bc_pe_992 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_992_clock),
    .reset(bc_pe_992_reset),
    .io_ho_input(bc_pe_992_io_ho_input),
    .io_ve_input(bc_pe_992_io_ve_input),
    .io_input_valid(bc_pe_992_io_input_valid),
    .io_iormac(bc_pe_992_io_iormac),
    .io_ve_out(bc_pe_992_io_ve_out),
    .io_ho_out(bc_pe_992_io_ho_out),
    .io_res_out(bc_pe_992_io_res_out)
  );
  bc_pe bc_pe_993 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_993_clock),
    .reset(bc_pe_993_reset),
    .io_ho_input(bc_pe_993_io_ho_input),
    .io_ve_input(bc_pe_993_io_ve_input),
    .io_input_valid(bc_pe_993_io_input_valid),
    .io_iormac(bc_pe_993_io_iormac),
    .io_ve_out(bc_pe_993_io_ve_out),
    .io_ho_out(bc_pe_993_io_ho_out),
    .io_res_out(bc_pe_993_io_res_out)
  );
  bc_pe bc_pe_994 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_994_clock),
    .reset(bc_pe_994_reset),
    .io_ho_input(bc_pe_994_io_ho_input),
    .io_ve_input(bc_pe_994_io_ve_input),
    .io_input_valid(bc_pe_994_io_input_valid),
    .io_iormac(bc_pe_994_io_iormac),
    .io_ve_out(bc_pe_994_io_ve_out),
    .io_ho_out(bc_pe_994_io_ho_out),
    .io_res_out(bc_pe_994_io_res_out)
  );
  bc_pe bc_pe_995 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_995_clock),
    .reset(bc_pe_995_reset),
    .io_ho_input(bc_pe_995_io_ho_input),
    .io_ve_input(bc_pe_995_io_ve_input),
    .io_input_valid(bc_pe_995_io_input_valid),
    .io_iormac(bc_pe_995_io_iormac),
    .io_ve_out(bc_pe_995_io_ve_out),
    .io_ho_out(bc_pe_995_io_ho_out),
    .io_res_out(bc_pe_995_io_res_out)
  );
  bc_pe bc_pe_996 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_996_clock),
    .reset(bc_pe_996_reset),
    .io_ho_input(bc_pe_996_io_ho_input),
    .io_ve_input(bc_pe_996_io_ve_input),
    .io_input_valid(bc_pe_996_io_input_valid),
    .io_iormac(bc_pe_996_io_iormac),
    .io_ve_out(bc_pe_996_io_ve_out),
    .io_ho_out(bc_pe_996_io_ho_out),
    .io_res_out(bc_pe_996_io_res_out)
  );
  bc_pe bc_pe_997 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_997_clock),
    .reset(bc_pe_997_reset),
    .io_ho_input(bc_pe_997_io_ho_input),
    .io_ve_input(bc_pe_997_io_ve_input),
    .io_input_valid(bc_pe_997_io_input_valid),
    .io_iormac(bc_pe_997_io_iormac),
    .io_ve_out(bc_pe_997_io_ve_out),
    .io_ho_out(bc_pe_997_io_ho_out),
    .io_res_out(bc_pe_997_io_res_out)
  );
  bc_pe bc_pe_998 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_998_clock),
    .reset(bc_pe_998_reset),
    .io_ho_input(bc_pe_998_io_ho_input),
    .io_ve_input(bc_pe_998_io_ve_input),
    .io_input_valid(bc_pe_998_io_input_valid),
    .io_iormac(bc_pe_998_io_iormac),
    .io_ve_out(bc_pe_998_io_ve_out),
    .io_ho_out(bc_pe_998_io_ho_out),
    .io_res_out(bc_pe_998_io_res_out)
  );
  bc_pe bc_pe_999 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_999_clock),
    .reset(bc_pe_999_reset),
    .io_ho_input(bc_pe_999_io_ho_input),
    .io_ve_input(bc_pe_999_io_ve_input),
    .io_input_valid(bc_pe_999_io_input_valid),
    .io_iormac(bc_pe_999_io_iormac),
    .io_ve_out(bc_pe_999_io_ve_out),
    .io_ho_out(bc_pe_999_io_ho_out),
    .io_res_out(bc_pe_999_io_res_out)
  );
  bc_pe bc_pe_1000 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1000_clock),
    .reset(bc_pe_1000_reset),
    .io_ho_input(bc_pe_1000_io_ho_input),
    .io_ve_input(bc_pe_1000_io_ve_input),
    .io_input_valid(bc_pe_1000_io_input_valid),
    .io_iormac(bc_pe_1000_io_iormac),
    .io_ve_out(bc_pe_1000_io_ve_out),
    .io_ho_out(bc_pe_1000_io_ho_out),
    .io_res_out(bc_pe_1000_io_res_out)
  );
  bc_pe bc_pe_1001 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1001_clock),
    .reset(bc_pe_1001_reset),
    .io_ho_input(bc_pe_1001_io_ho_input),
    .io_ve_input(bc_pe_1001_io_ve_input),
    .io_input_valid(bc_pe_1001_io_input_valid),
    .io_iormac(bc_pe_1001_io_iormac),
    .io_ve_out(bc_pe_1001_io_ve_out),
    .io_ho_out(bc_pe_1001_io_ho_out),
    .io_res_out(bc_pe_1001_io_res_out)
  );
  bc_pe bc_pe_1002 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1002_clock),
    .reset(bc_pe_1002_reset),
    .io_ho_input(bc_pe_1002_io_ho_input),
    .io_ve_input(bc_pe_1002_io_ve_input),
    .io_input_valid(bc_pe_1002_io_input_valid),
    .io_iormac(bc_pe_1002_io_iormac),
    .io_ve_out(bc_pe_1002_io_ve_out),
    .io_ho_out(bc_pe_1002_io_ho_out),
    .io_res_out(bc_pe_1002_io_res_out)
  );
  bc_pe bc_pe_1003 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1003_clock),
    .reset(bc_pe_1003_reset),
    .io_ho_input(bc_pe_1003_io_ho_input),
    .io_ve_input(bc_pe_1003_io_ve_input),
    .io_input_valid(bc_pe_1003_io_input_valid),
    .io_iormac(bc_pe_1003_io_iormac),
    .io_ve_out(bc_pe_1003_io_ve_out),
    .io_ho_out(bc_pe_1003_io_ho_out),
    .io_res_out(bc_pe_1003_io_res_out)
  );
  bc_pe bc_pe_1004 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1004_clock),
    .reset(bc_pe_1004_reset),
    .io_ho_input(bc_pe_1004_io_ho_input),
    .io_ve_input(bc_pe_1004_io_ve_input),
    .io_input_valid(bc_pe_1004_io_input_valid),
    .io_iormac(bc_pe_1004_io_iormac),
    .io_ve_out(bc_pe_1004_io_ve_out),
    .io_ho_out(bc_pe_1004_io_ho_out),
    .io_res_out(bc_pe_1004_io_res_out)
  );
  bc_pe bc_pe_1005 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1005_clock),
    .reset(bc_pe_1005_reset),
    .io_ho_input(bc_pe_1005_io_ho_input),
    .io_ve_input(bc_pe_1005_io_ve_input),
    .io_input_valid(bc_pe_1005_io_input_valid),
    .io_iormac(bc_pe_1005_io_iormac),
    .io_ve_out(bc_pe_1005_io_ve_out),
    .io_ho_out(bc_pe_1005_io_ho_out),
    .io_res_out(bc_pe_1005_io_res_out)
  );
  bc_pe bc_pe_1006 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1006_clock),
    .reset(bc_pe_1006_reset),
    .io_ho_input(bc_pe_1006_io_ho_input),
    .io_ve_input(bc_pe_1006_io_ve_input),
    .io_input_valid(bc_pe_1006_io_input_valid),
    .io_iormac(bc_pe_1006_io_iormac),
    .io_ve_out(bc_pe_1006_io_ve_out),
    .io_ho_out(bc_pe_1006_io_ho_out),
    .io_res_out(bc_pe_1006_io_res_out)
  );
  bc_pe bc_pe_1007 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1007_clock),
    .reset(bc_pe_1007_reset),
    .io_ho_input(bc_pe_1007_io_ho_input),
    .io_ve_input(bc_pe_1007_io_ve_input),
    .io_input_valid(bc_pe_1007_io_input_valid),
    .io_iormac(bc_pe_1007_io_iormac),
    .io_ve_out(bc_pe_1007_io_ve_out),
    .io_ho_out(bc_pe_1007_io_ho_out),
    .io_res_out(bc_pe_1007_io_res_out)
  );
  bc_pe bc_pe_1008 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1008_clock),
    .reset(bc_pe_1008_reset),
    .io_ho_input(bc_pe_1008_io_ho_input),
    .io_ve_input(bc_pe_1008_io_ve_input),
    .io_input_valid(bc_pe_1008_io_input_valid),
    .io_iormac(bc_pe_1008_io_iormac),
    .io_ve_out(bc_pe_1008_io_ve_out),
    .io_ho_out(bc_pe_1008_io_ho_out),
    .io_res_out(bc_pe_1008_io_res_out)
  );
  bc_pe bc_pe_1009 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1009_clock),
    .reset(bc_pe_1009_reset),
    .io_ho_input(bc_pe_1009_io_ho_input),
    .io_ve_input(bc_pe_1009_io_ve_input),
    .io_input_valid(bc_pe_1009_io_input_valid),
    .io_iormac(bc_pe_1009_io_iormac),
    .io_ve_out(bc_pe_1009_io_ve_out),
    .io_ho_out(bc_pe_1009_io_ho_out),
    .io_res_out(bc_pe_1009_io_res_out)
  );
  bc_pe bc_pe_1010 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1010_clock),
    .reset(bc_pe_1010_reset),
    .io_ho_input(bc_pe_1010_io_ho_input),
    .io_ve_input(bc_pe_1010_io_ve_input),
    .io_input_valid(bc_pe_1010_io_input_valid),
    .io_iormac(bc_pe_1010_io_iormac),
    .io_ve_out(bc_pe_1010_io_ve_out),
    .io_ho_out(bc_pe_1010_io_ho_out),
    .io_res_out(bc_pe_1010_io_res_out)
  );
  bc_pe bc_pe_1011 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1011_clock),
    .reset(bc_pe_1011_reset),
    .io_ho_input(bc_pe_1011_io_ho_input),
    .io_ve_input(bc_pe_1011_io_ve_input),
    .io_input_valid(bc_pe_1011_io_input_valid),
    .io_iormac(bc_pe_1011_io_iormac),
    .io_ve_out(bc_pe_1011_io_ve_out),
    .io_ho_out(bc_pe_1011_io_ho_out),
    .io_res_out(bc_pe_1011_io_res_out)
  );
  bc_pe bc_pe_1012 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1012_clock),
    .reset(bc_pe_1012_reset),
    .io_ho_input(bc_pe_1012_io_ho_input),
    .io_ve_input(bc_pe_1012_io_ve_input),
    .io_input_valid(bc_pe_1012_io_input_valid),
    .io_iormac(bc_pe_1012_io_iormac),
    .io_ve_out(bc_pe_1012_io_ve_out),
    .io_ho_out(bc_pe_1012_io_ho_out),
    .io_res_out(bc_pe_1012_io_res_out)
  );
  bc_pe bc_pe_1013 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1013_clock),
    .reset(bc_pe_1013_reset),
    .io_ho_input(bc_pe_1013_io_ho_input),
    .io_ve_input(bc_pe_1013_io_ve_input),
    .io_input_valid(bc_pe_1013_io_input_valid),
    .io_iormac(bc_pe_1013_io_iormac),
    .io_ve_out(bc_pe_1013_io_ve_out),
    .io_ho_out(bc_pe_1013_io_ho_out),
    .io_res_out(bc_pe_1013_io_res_out)
  );
  bc_pe bc_pe_1014 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1014_clock),
    .reset(bc_pe_1014_reset),
    .io_ho_input(bc_pe_1014_io_ho_input),
    .io_ve_input(bc_pe_1014_io_ve_input),
    .io_input_valid(bc_pe_1014_io_input_valid),
    .io_iormac(bc_pe_1014_io_iormac),
    .io_ve_out(bc_pe_1014_io_ve_out),
    .io_ho_out(bc_pe_1014_io_ho_out),
    .io_res_out(bc_pe_1014_io_res_out)
  );
  bc_pe bc_pe_1015 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1015_clock),
    .reset(bc_pe_1015_reset),
    .io_ho_input(bc_pe_1015_io_ho_input),
    .io_ve_input(bc_pe_1015_io_ve_input),
    .io_input_valid(bc_pe_1015_io_input_valid),
    .io_iormac(bc_pe_1015_io_iormac),
    .io_ve_out(bc_pe_1015_io_ve_out),
    .io_ho_out(bc_pe_1015_io_ho_out),
    .io_res_out(bc_pe_1015_io_res_out)
  );
  bc_pe bc_pe_1016 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1016_clock),
    .reset(bc_pe_1016_reset),
    .io_ho_input(bc_pe_1016_io_ho_input),
    .io_ve_input(bc_pe_1016_io_ve_input),
    .io_input_valid(bc_pe_1016_io_input_valid),
    .io_iormac(bc_pe_1016_io_iormac),
    .io_ve_out(bc_pe_1016_io_ve_out),
    .io_ho_out(bc_pe_1016_io_ho_out),
    .io_res_out(bc_pe_1016_io_res_out)
  );
  bc_pe bc_pe_1017 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1017_clock),
    .reset(bc_pe_1017_reset),
    .io_ho_input(bc_pe_1017_io_ho_input),
    .io_ve_input(bc_pe_1017_io_ve_input),
    .io_input_valid(bc_pe_1017_io_input_valid),
    .io_iormac(bc_pe_1017_io_iormac),
    .io_ve_out(bc_pe_1017_io_ve_out),
    .io_ho_out(bc_pe_1017_io_ho_out),
    .io_res_out(bc_pe_1017_io_res_out)
  );
  bc_pe bc_pe_1018 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1018_clock),
    .reset(bc_pe_1018_reset),
    .io_ho_input(bc_pe_1018_io_ho_input),
    .io_ve_input(bc_pe_1018_io_ve_input),
    .io_input_valid(bc_pe_1018_io_input_valid),
    .io_iormac(bc_pe_1018_io_iormac),
    .io_ve_out(bc_pe_1018_io_ve_out),
    .io_ho_out(bc_pe_1018_io_ho_out),
    .io_res_out(bc_pe_1018_io_res_out)
  );
  bc_pe bc_pe_1019 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1019_clock),
    .reset(bc_pe_1019_reset),
    .io_ho_input(bc_pe_1019_io_ho_input),
    .io_ve_input(bc_pe_1019_io_ve_input),
    .io_input_valid(bc_pe_1019_io_input_valid),
    .io_iormac(bc_pe_1019_io_iormac),
    .io_ve_out(bc_pe_1019_io_ve_out),
    .io_ho_out(bc_pe_1019_io_ho_out),
    .io_res_out(bc_pe_1019_io_res_out)
  );
  bc_pe bc_pe_1020 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1020_clock),
    .reset(bc_pe_1020_reset),
    .io_ho_input(bc_pe_1020_io_ho_input),
    .io_ve_input(bc_pe_1020_io_ve_input),
    .io_input_valid(bc_pe_1020_io_input_valid),
    .io_iormac(bc_pe_1020_io_iormac),
    .io_ve_out(bc_pe_1020_io_ve_out),
    .io_ho_out(bc_pe_1020_io_ho_out),
    .io_res_out(bc_pe_1020_io_res_out)
  );
  bc_pe bc_pe_1021 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1021_clock),
    .reset(bc_pe_1021_reset),
    .io_ho_input(bc_pe_1021_io_ho_input),
    .io_ve_input(bc_pe_1021_io_ve_input),
    .io_input_valid(bc_pe_1021_io_input_valid),
    .io_iormac(bc_pe_1021_io_iormac),
    .io_ve_out(bc_pe_1021_io_ve_out),
    .io_ho_out(bc_pe_1021_io_ho_out),
    .io_res_out(bc_pe_1021_io_res_out)
  );
  bc_pe bc_pe_1022 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1022_clock),
    .reset(bc_pe_1022_reset),
    .io_ho_input(bc_pe_1022_io_ho_input),
    .io_ve_input(bc_pe_1022_io_ve_input),
    .io_input_valid(bc_pe_1022_io_input_valid),
    .io_iormac(bc_pe_1022_io_iormac),
    .io_ve_out(bc_pe_1022_io_ve_out),
    .io_ho_out(bc_pe_1022_io_ho_out),
    .io_res_out(bc_pe_1022_io_res_out)
  );
  bc_pe bc_pe_1023 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1023_clock),
    .reset(bc_pe_1023_reset),
    .io_ho_input(bc_pe_1023_io_ho_input),
    .io_ve_input(bc_pe_1023_io_ve_input),
    .io_input_valid(bc_pe_1023_io_input_valid),
    .io_iormac(bc_pe_1023_io_iormac),
    .io_ve_out(bc_pe_1023_io_ve_out),
    .io_ho_out(bc_pe_1023_io_ho_out),
    .io_res_out(bc_pe_1023_io_res_out)
  );
  assign io_out_0 = bc_pe_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1 = bc_pe_1_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_2 = bc_pe_2_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_3 = bc_pe_3_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_4 = bc_pe_4_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_5 = bc_pe_5_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_6 = bc_pe_6_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_7 = bc_pe_7_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_8 = bc_pe_8_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_9 = bc_pe_9_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_10 = bc_pe_10_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_11 = bc_pe_11_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_12 = bc_pe_12_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_13 = bc_pe_13_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_14 = bc_pe_14_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_15 = bc_pe_15_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_16 = bc_pe_16_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_17 = bc_pe_17_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_18 = bc_pe_18_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_19 = bc_pe_19_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_20 = bc_pe_20_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_21 = bc_pe_21_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_22 = bc_pe_22_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_23 = bc_pe_23_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_24 = bc_pe_24_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_25 = bc_pe_25_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_26 = bc_pe_26_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_27 = bc_pe_27_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_28 = bc_pe_28_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_29 = bc_pe_29_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_30 = bc_pe_30_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_31 = bc_pe_31_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_32 = bc_pe_32_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_33 = bc_pe_33_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_34 = bc_pe_34_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_35 = bc_pe_35_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_36 = bc_pe_36_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_37 = bc_pe_37_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_38 = bc_pe_38_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_39 = bc_pe_39_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_40 = bc_pe_40_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_41 = bc_pe_41_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_42 = bc_pe_42_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_43 = bc_pe_43_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_44 = bc_pe_44_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_45 = bc_pe_45_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_46 = bc_pe_46_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_47 = bc_pe_47_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_48 = bc_pe_48_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_49 = bc_pe_49_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_50 = bc_pe_50_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_51 = bc_pe_51_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_52 = bc_pe_52_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_53 = bc_pe_53_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_54 = bc_pe_54_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_55 = bc_pe_55_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_56 = bc_pe_56_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_57 = bc_pe_57_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_58 = bc_pe_58_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_59 = bc_pe_59_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_60 = bc_pe_60_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_61 = bc_pe_61_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_62 = bc_pe_62_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_63 = bc_pe_63_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_64 = bc_pe_64_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_65 = bc_pe_65_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_66 = bc_pe_66_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_67 = bc_pe_67_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_68 = bc_pe_68_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_69 = bc_pe_69_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_70 = bc_pe_70_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_71 = bc_pe_71_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_72 = bc_pe_72_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_73 = bc_pe_73_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_74 = bc_pe_74_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_75 = bc_pe_75_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_76 = bc_pe_76_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_77 = bc_pe_77_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_78 = bc_pe_78_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_79 = bc_pe_79_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_80 = bc_pe_80_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_81 = bc_pe_81_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_82 = bc_pe_82_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_83 = bc_pe_83_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_84 = bc_pe_84_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_85 = bc_pe_85_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_86 = bc_pe_86_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_87 = bc_pe_87_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_88 = bc_pe_88_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_89 = bc_pe_89_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_90 = bc_pe_90_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_91 = bc_pe_91_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_92 = bc_pe_92_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_93 = bc_pe_93_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_94 = bc_pe_94_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_95 = bc_pe_95_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_96 = bc_pe_96_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_97 = bc_pe_97_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_98 = bc_pe_98_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_99 = bc_pe_99_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_100 = bc_pe_100_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_101 = bc_pe_101_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_102 = bc_pe_102_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_103 = bc_pe_103_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_104 = bc_pe_104_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_105 = bc_pe_105_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_106 = bc_pe_106_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_107 = bc_pe_107_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_108 = bc_pe_108_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_109 = bc_pe_109_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_110 = bc_pe_110_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_111 = bc_pe_111_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_112 = bc_pe_112_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_113 = bc_pe_113_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_114 = bc_pe_114_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_115 = bc_pe_115_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_116 = bc_pe_116_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_117 = bc_pe_117_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_118 = bc_pe_118_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_119 = bc_pe_119_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_120 = bc_pe_120_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_121 = bc_pe_121_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_122 = bc_pe_122_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_123 = bc_pe_123_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_124 = bc_pe_124_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_125 = bc_pe_125_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_126 = bc_pe_126_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_127 = bc_pe_127_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_128 = bc_pe_128_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_129 = bc_pe_129_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_130 = bc_pe_130_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_131 = bc_pe_131_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_132 = bc_pe_132_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_133 = bc_pe_133_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_134 = bc_pe_134_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_135 = bc_pe_135_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_136 = bc_pe_136_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_137 = bc_pe_137_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_138 = bc_pe_138_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_139 = bc_pe_139_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_140 = bc_pe_140_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_141 = bc_pe_141_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_142 = bc_pe_142_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_143 = bc_pe_143_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_144 = bc_pe_144_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_145 = bc_pe_145_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_146 = bc_pe_146_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_147 = bc_pe_147_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_148 = bc_pe_148_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_149 = bc_pe_149_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_150 = bc_pe_150_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_151 = bc_pe_151_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_152 = bc_pe_152_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_153 = bc_pe_153_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_154 = bc_pe_154_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_155 = bc_pe_155_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_156 = bc_pe_156_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_157 = bc_pe_157_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_158 = bc_pe_158_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_159 = bc_pe_159_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_160 = bc_pe_160_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_161 = bc_pe_161_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_162 = bc_pe_162_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_163 = bc_pe_163_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_164 = bc_pe_164_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_165 = bc_pe_165_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_166 = bc_pe_166_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_167 = bc_pe_167_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_168 = bc_pe_168_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_169 = bc_pe_169_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_170 = bc_pe_170_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_171 = bc_pe_171_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_172 = bc_pe_172_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_173 = bc_pe_173_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_174 = bc_pe_174_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_175 = bc_pe_175_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_176 = bc_pe_176_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_177 = bc_pe_177_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_178 = bc_pe_178_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_179 = bc_pe_179_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_180 = bc_pe_180_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_181 = bc_pe_181_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_182 = bc_pe_182_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_183 = bc_pe_183_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_184 = bc_pe_184_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_185 = bc_pe_185_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_186 = bc_pe_186_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_187 = bc_pe_187_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_188 = bc_pe_188_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_189 = bc_pe_189_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_190 = bc_pe_190_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_191 = bc_pe_191_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_192 = bc_pe_192_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_193 = bc_pe_193_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_194 = bc_pe_194_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_195 = bc_pe_195_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_196 = bc_pe_196_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_197 = bc_pe_197_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_198 = bc_pe_198_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_199 = bc_pe_199_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_200 = bc_pe_200_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_201 = bc_pe_201_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_202 = bc_pe_202_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_203 = bc_pe_203_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_204 = bc_pe_204_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_205 = bc_pe_205_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_206 = bc_pe_206_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_207 = bc_pe_207_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_208 = bc_pe_208_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_209 = bc_pe_209_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_210 = bc_pe_210_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_211 = bc_pe_211_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_212 = bc_pe_212_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_213 = bc_pe_213_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_214 = bc_pe_214_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_215 = bc_pe_215_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_216 = bc_pe_216_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_217 = bc_pe_217_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_218 = bc_pe_218_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_219 = bc_pe_219_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_220 = bc_pe_220_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_221 = bc_pe_221_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_222 = bc_pe_222_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_223 = bc_pe_223_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_224 = bc_pe_224_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_225 = bc_pe_225_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_226 = bc_pe_226_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_227 = bc_pe_227_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_228 = bc_pe_228_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_229 = bc_pe_229_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_230 = bc_pe_230_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_231 = bc_pe_231_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_232 = bc_pe_232_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_233 = bc_pe_233_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_234 = bc_pe_234_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_235 = bc_pe_235_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_236 = bc_pe_236_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_237 = bc_pe_237_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_238 = bc_pe_238_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_239 = bc_pe_239_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_240 = bc_pe_240_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_241 = bc_pe_241_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_242 = bc_pe_242_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_243 = bc_pe_243_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_244 = bc_pe_244_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_245 = bc_pe_245_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_246 = bc_pe_246_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_247 = bc_pe_247_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_248 = bc_pe_248_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_249 = bc_pe_249_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_250 = bc_pe_250_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_251 = bc_pe_251_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_252 = bc_pe_252_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_253 = bc_pe_253_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_254 = bc_pe_254_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_255 = bc_pe_255_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_256 = bc_pe_256_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_257 = bc_pe_257_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_258 = bc_pe_258_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_259 = bc_pe_259_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_260 = bc_pe_260_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_261 = bc_pe_261_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_262 = bc_pe_262_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_263 = bc_pe_263_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_264 = bc_pe_264_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_265 = bc_pe_265_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_266 = bc_pe_266_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_267 = bc_pe_267_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_268 = bc_pe_268_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_269 = bc_pe_269_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_270 = bc_pe_270_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_271 = bc_pe_271_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_272 = bc_pe_272_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_273 = bc_pe_273_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_274 = bc_pe_274_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_275 = bc_pe_275_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_276 = bc_pe_276_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_277 = bc_pe_277_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_278 = bc_pe_278_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_279 = bc_pe_279_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_280 = bc_pe_280_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_281 = bc_pe_281_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_282 = bc_pe_282_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_283 = bc_pe_283_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_284 = bc_pe_284_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_285 = bc_pe_285_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_286 = bc_pe_286_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_287 = bc_pe_287_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_288 = bc_pe_288_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_289 = bc_pe_289_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_290 = bc_pe_290_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_291 = bc_pe_291_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_292 = bc_pe_292_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_293 = bc_pe_293_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_294 = bc_pe_294_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_295 = bc_pe_295_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_296 = bc_pe_296_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_297 = bc_pe_297_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_298 = bc_pe_298_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_299 = bc_pe_299_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_300 = bc_pe_300_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_301 = bc_pe_301_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_302 = bc_pe_302_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_303 = bc_pe_303_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_304 = bc_pe_304_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_305 = bc_pe_305_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_306 = bc_pe_306_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_307 = bc_pe_307_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_308 = bc_pe_308_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_309 = bc_pe_309_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_310 = bc_pe_310_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_311 = bc_pe_311_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_312 = bc_pe_312_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_313 = bc_pe_313_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_314 = bc_pe_314_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_315 = bc_pe_315_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_316 = bc_pe_316_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_317 = bc_pe_317_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_318 = bc_pe_318_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_319 = bc_pe_319_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_320 = bc_pe_320_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_321 = bc_pe_321_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_322 = bc_pe_322_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_323 = bc_pe_323_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_324 = bc_pe_324_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_325 = bc_pe_325_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_326 = bc_pe_326_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_327 = bc_pe_327_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_328 = bc_pe_328_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_329 = bc_pe_329_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_330 = bc_pe_330_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_331 = bc_pe_331_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_332 = bc_pe_332_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_333 = bc_pe_333_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_334 = bc_pe_334_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_335 = bc_pe_335_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_336 = bc_pe_336_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_337 = bc_pe_337_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_338 = bc_pe_338_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_339 = bc_pe_339_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_340 = bc_pe_340_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_341 = bc_pe_341_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_342 = bc_pe_342_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_343 = bc_pe_343_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_344 = bc_pe_344_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_345 = bc_pe_345_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_346 = bc_pe_346_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_347 = bc_pe_347_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_348 = bc_pe_348_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_349 = bc_pe_349_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_350 = bc_pe_350_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_351 = bc_pe_351_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_352 = bc_pe_352_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_353 = bc_pe_353_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_354 = bc_pe_354_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_355 = bc_pe_355_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_356 = bc_pe_356_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_357 = bc_pe_357_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_358 = bc_pe_358_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_359 = bc_pe_359_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_360 = bc_pe_360_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_361 = bc_pe_361_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_362 = bc_pe_362_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_363 = bc_pe_363_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_364 = bc_pe_364_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_365 = bc_pe_365_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_366 = bc_pe_366_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_367 = bc_pe_367_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_368 = bc_pe_368_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_369 = bc_pe_369_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_370 = bc_pe_370_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_371 = bc_pe_371_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_372 = bc_pe_372_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_373 = bc_pe_373_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_374 = bc_pe_374_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_375 = bc_pe_375_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_376 = bc_pe_376_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_377 = bc_pe_377_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_378 = bc_pe_378_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_379 = bc_pe_379_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_380 = bc_pe_380_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_381 = bc_pe_381_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_382 = bc_pe_382_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_383 = bc_pe_383_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_384 = bc_pe_384_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_385 = bc_pe_385_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_386 = bc_pe_386_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_387 = bc_pe_387_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_388 = bc_pe_388_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_389 = bc_pe_389_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_390 = bc_pe_390_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_391 = bc_pe_391_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_392 = bc_pe_392_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_393 = bc_pe_393_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_394 = bc_pe_394_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_395 = bc_pe_395_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_396 = bc_pe_396_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_397 = bc_pe_397_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_398 = bc_pe_398_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_399 = bc_pe_399_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_400 = bc_pe_400_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_401 = bc_pe_401_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_402 = bc_pe_402_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_403 = bc_pe_403_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_404 = bc_pe_404_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_405 = bc_pe_405_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_406 = bc_pe_406_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_407 = bc_pe_407_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_408 = bc_pe_408_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_409 = bc_pe_409_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_410 = bc_pe_410_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_411 = bc_pe_411_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_412 = bc_pe_412_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_413 = bc_pe_413_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_414 = bc_pe_414_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_415 = bc_pe_415_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_416 = bc_pe_416_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_417 = bc_pe_417_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_418 = bc_pe_418_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_419 = bc_pe_419_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_420 = bc_pe_420_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_421 = bc_pe_421_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_422 = bc_pe_422_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_423 = bc_pe_423_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_424 = bc_pe_424_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_425 = bc_pe_425_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_426 = bc_pe_426_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_427 = bc_pe_427_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_428 = bc_pe_428_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_429 = bc_pe_429_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_430 = bc_pe_430_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_431 = bc_pe_431_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_432 = bc_pe_432_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_433 = bc_pe_433_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_434 = bc_pe_434_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_435 = bc_pe_435_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_436 = bc_pe_436_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_437 = bc_pe_437_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_438 = bc_pe_438_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_439 = bc_pe_439_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_440 = bc_pe_440_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_441 = bc_pe_441_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_442 = bc_pe_442_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_443 = bc_pe_443_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_444 = bc_pe_444_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_445 = bc_pe_445_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_446 = bc_pe_446_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_447 = bc_pe_447_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_448 = bc_pe_448_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_449 = bc_pe_449_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_450 = bc_pe_450_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_451 = bc_pe_451_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_452 = bc_pe_452_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_453 = bc_pe_453_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_454 = bc_pe_454_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_455 = bc_pe_455_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_456 = bc_pe_456_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_457 = bc_pe_457_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_458 = bc_pe_458_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_459 = bc_pe_459_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_460 = bc_pe_460_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_461 = bc_pe_461_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_462 = bc_pe_462_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_463 = bc_pe_463_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_464 = bc_pe_464_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_465 = bc_pe_465_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_466 = bc_pe_466_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_467 = bc_pe_467_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_468 = bc_pe_468_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_469 = bc_pe_469_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_470 = bc_pe_470_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_471 = bc_pe_471_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_472 = bc_pe_472_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_473 = bc_pe_473_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_474 = bc_pe_474_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_475 = bc_pe_475_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_476 = bc_pe_476_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_477 = bc_pe_477_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_478 = bc_pe_478_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_479 = bc_pe_479_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_480 = bc_pe_480_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_481 = bc_pe_481_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_482 = bc_pe_482_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_483 = bc_pe_483_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_484 = bc_pe_484_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_485 = bc_pe_485_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_486 = bc_pe_486_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_487 = bc_pe_487_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_488 = bc_pe_488_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_489 = bc_pe_489_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_490 = bc_pe_490_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_491 = bc_pe_491_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_492 = bc_pe_492_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_493 = bc_pe_493_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_494 = bc_pe_494_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_495 = bc_pe_495_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_496 = bc_pe_496_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_497 = bc_pe_497_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_498 = bc_pe_498_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_499 = bc_pe_499_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_500 = bc_pe_500_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_501 = bc_pe_501_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_502 = bc_pe_502_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_503 = bc_pe_503_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_504 = bc_pe_504_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_505 = bc_pe_505_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_506 = bc_pe_506_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_507 = bc_pe_507_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_508 = bc_pe_508_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_509 = bc_pe_509_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_510 = bc_pe_510_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_511 = bc_pe_511_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_512 = bc_pe_512_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_513 = bc_pe_513_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_514 = bc_pe_514_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_515 = bc_pe_515_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_516 = bc_pe_516_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_517 = bc_pe_517_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_518 = bc_pe_518_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_519 = bc_pe_519_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_520 = bc_pe_520_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_521 = bc_pe_521_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_522 = bc_pe_522_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_523 = bc_pe_523_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_524 = bc_pe_524_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_525 = bc_pe_525_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_526 = bc_pe_526_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_527 = bc_pe_527_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_528 = bc_pe_528_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_529 = bc_pe_529_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_530 = bc_pe_530_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_531 = bc_pe_531_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_532 = bc_pe_532_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_533 = bc_pe_533_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_534 = bc_pe_534_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_535 = bc_pe_535_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_536 = bc_pe_536_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_537 = bc_pe_537_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_538 = bc_pe_538_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_539 = bc_pe_539_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_540 = bc_pe_540_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_541 = bc_pe_541_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_542 = bc_pe_542_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_543 = bc_pe_543_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_544 = bc_pe_544_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_545 = bc_pe_545_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_546 = bc_pe_546_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_547 = bc_pe_547_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_548 = bc_pe_548_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_549 = bc_pe_549_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_550 = bc_pe_550_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_551 = bc_pe_551_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_552 = bc_pe_552_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_553 = bc_pe_553_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_554 = bc_pe_554_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_555 = bc_pe_555_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_556 = bc_pe_556_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_557 = bc_pe_557_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_558 = bc_pe_558_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_559 = bc_pe_559_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_560 = bc_pe_560_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_561 = bc_pe_561_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_562 = bc_pe_562_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_563 = bc_pe_563_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_564 = bc_pe_564_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_565 = bc_pe_565_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_566 = bc_pe_566_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_567 = bc_pe_567_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_568 = bc_pe_568_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_569 = bc_pe_569_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_570 = bc_pe_570_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_571 = bc_pe_571_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_572 = bc_pe_572_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_573 = bc_pe_573_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_574 = bc_pe_574_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_575 = bc_pe_575_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_576 = bc_pe_576_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_577 = bc_pe_577_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_578 = bc_pe_578_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_579 = bc_pe_579_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_580 = bc_pe_580_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_581 = bc_pe_581_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_582 = bc_pe_582_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_583 = bc_pe_583_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_584 = bc_pe_584_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_585 = bc_pe_585_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_586 = bc_pe_586_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_587 = bc_pe_587_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_588 = bc_pe_588_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_589 = bc_pe_589_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_590 = bc_pe_590_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_591 = bc_pe_591_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_592 = bc_pe_592_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_593 = bc_pe_593_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_594 = bc_pe_594_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_595 = bc_pe_595_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_596 = bc_pe_596_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_597 = bc_pe_597_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_598 = bc_pe_598_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_599 = bc_pe_599_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_600 = bc_pe_600_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_601 = bc_pe_601_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_602 = bc_pe_602_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_603 = bc_pe_603_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_604 = bc_pe_604_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_605 = bc_pe_605_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_606 = bc_pe_606_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_607 = bc_pe_607_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_608 = bc_pe_608_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_609 = bc_pe_609_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_610 = bc_pe_610_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_611 = bc_pe_611_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_612 = bc_pe_612_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_613 = bc_pe_613_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_614 = bc_pe_614_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_615 = bc_pe_615_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_616 = bc_pe_616_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_617 = bc_pe_617_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_618 = bc_pe_618_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_619 = bc_pe_619_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_620 = bc_pe_620_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_621 = bc_pe_621_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_622 = bc_pe_622_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_623 = bc_pe_623_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_624 = bc_pe_624_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_625 = bc_pe_625_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_626 = bc_pe_626_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_627 = bc_pe_627_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_628 = bc_pe_628_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_629 = bc_pe_629_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_630 = bc_pe_630_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_631 = bc_pe_631_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_632 = bc_pe_632_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_633 = bc_pe_633_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_634 = bc_pe_634_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_635 = bc_pe_635_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_636 = bc_pe_636_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_637 = bc_pe_637_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_638 = bc_pe_638_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_639 = bc_pe_639_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_640 = bc_pe_640_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_641 = bc_pe_641_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_642 = bc_pe_642_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_643 = bc_pe_643_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_644 = bc_pe_644_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_645 = bc_pe_645_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_646 = bc_pe_646_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_647 = bc_pe_647_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_648 = bc_pe_648_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_649 = bc_pe_649_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_650 = bc_pe_650_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_651 = bc_pe_651_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_652 = bc_pe_652_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_653 = bc_pe_653_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_654 = bc_pe_654_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_655 = bc_pe_655_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_656 = bc_pe_656_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_657 = bc_pe_657_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_658 = bc_pe_658_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_659 = bc_pe_659_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_660 = bc_pe_660_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_661 = bc_pe_661_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_662 = bc_pe_662_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_663 = bc_pe_663_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_664 = bc_pe_664_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_665 = bc_pe_665_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_666 = bc_pe_666_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_667 = bc_pe_667_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_668 = bc_pe_668_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_669 = bc_pe_669_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_670 = bc_pe_670_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_671 = bc_pe_671_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_672 = bc_pe_672_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_673 = bc_pe_673_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_674 = bc_pe_674_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_675 = bc_pe_675_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_676 = bc_pe_676_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_677 = bc_pe_677_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_678 = bc_pe_678_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_679 = bc_pe_679_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_680 = bc_pe_680_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_681 = bc_pe_681_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_682 = bc_pe_682_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_683 = bc_pe_683_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_684 = bc_pe_684_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_685 = bc_pe_685_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_686 = bc_pe_686_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_687 = bc_pe_687_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_688 = bc_pe_688_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_689 = bc_pe_689_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_690 = bc_pe_690_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_691 = bc_pe_691_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_692 = bc_pe_692_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_693 = bc_pe_693_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_694 = bc_pe_694_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_695 = bc_pe_695_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_696 = bc_pe_696_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_697 = bc_pe_697_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_698 = bc_pe_698_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_699 = bc_pe_699_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_700 = bc_pe_700_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_701 = bc_pe_701_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_702 = bc_pe_702_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_703 = bc_pe_703_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_704 = bc_pe_704_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_705 = bc_pe_705_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_706 = bc_pe_706_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_707 = bc_pe_707_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_708 = bc_pe_708_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_709 = bc_pe_709_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_710 = bc_pe_710_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_711 = bc_pe_711_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_712 = bc_pe_712_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_713 = bc_pe_713_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_714 = bc_pe_714_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_715 = bc_pe_715_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_716 = bc_pe_716_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_717 = bc_pe_717_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_718 = bc_pe_718_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_719 = bc_pe_719_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_720 = bc_pe_720_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_721 = bc_pe_721_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_722 = bc_pe_722_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_723 = bc_pe_723_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_724 = bc_pe_724_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_725 = bc_pe_725_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_726 = bc_pe_726_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_727 = bc_pe_727_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_728 = bc_pe_728_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_729 = bc_pe_729_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_730 = bc_pe_730_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_731 = bc_pe_731_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_732 = bc_pe_732_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_733 = bc_pe_733_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_734 = bc_pe_734_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_735 = bc_pe_735_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_736 = bc_pe_736_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_737 = bc_pe_737_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_738 = bc_pe_738_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_739 = bc_pe_739_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_740 = bc_pe_740_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_741 = bc_pe_741_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_742 = bc_pe_742_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_743 = bc_pe_743_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_744 = bc_pe_744_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_745 = bc_pe_745_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_746 = bc_pe_746_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_747 = bc_pe_747_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_748 = bc_pe_748_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_749 = bc_pe_749_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_750 = bc_pe_750_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_751 = bc_pe_751_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_752 = bc_pe_752_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_753 = bc_pe_753_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_754 = bc_pe_754_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_755 = bc_pe_755_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_756 = bc_pe_756_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_757 = bc_pe_757_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_758 = bc_pe_758_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_759 = bc_pe_759_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_760 = bc_pe_760_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_761 = bc_pe_761_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_762 = bc_pe_762_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_763 = bc_pe_763_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_764 = bc_pe_764_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_765 = bc_pe_765_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_766 = bc_pe_766_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_767 = bc_pe_767_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_768 = bc_pe_768_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_769 = bc_pe_769_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_770 = bc_pe_770_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_771 = bc_pe_771_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_772 = bc_pe_772_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_773 = bc_pe_773_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_774 = bc_pe_774_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_775 = bc_pe_775_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_776 = bc_pe_776_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_777 = bc_pe_777_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_778 = bc_pe_778_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_779 = bc_pe_779_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_780 = bc_pe_780_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_781 = bc_pe_781_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_782 = bc_pe_782_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_783 = bc_pe_783_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_784 = bc_pe_784_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_785 = bc_pe_785_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_786 = bc_pe_786_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_787 = bc_pe_787_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_788 = bc_pe_788_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_789 = bc_pe_789_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_790 = bc_pe_790_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_791 = bc_pe_791_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_792 = bc_pe_792_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_793 = bc_pe_793_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_794 = bc_pe_794_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_795 = bc_pe_795_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_796 = bc_pe_796_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_797 = bc_pe_797_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_798 = bc_pe_798_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_799 = bc_pe_799_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_800 = bc_pe_800_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_801 = bc_pe_801_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_802 = bc_pe_802_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_803 = bc_pe_803_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_804 = bc_pe_804_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_805 = bc_pe_805_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_806 = bc_pe_806_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_807 = bc_pe_807_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_808 = bc_pe_808_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_809 = bc_pe_809_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_810 = bc_pe_810_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_811 = bc_pe_811_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_812 = bc_pe_812_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_813 = bc_pe_813_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_814 = bc_pe_814_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_815 = bc_pe_815_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_816 = bc_pe_816_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_817 = bc_pe_817_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_818 = bc_pe_818_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_819 = bc_pe_819_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_820 = bc_pe_820_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_821 = bc_pe_821_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_822 = bc_pe_822_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_823 = bc_pe_823_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_824 = bc_pe_824_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_825 = bc_pe_825_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_826 = bc_pe_826_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_827 = bc_pe_827_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_828 = bc_pe_828_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_829 = bc_pe_829_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_830 = bc_pe_830_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_831 = bc_pe_831_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_832 = bc_pe_832_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_833 = bc_pe_833_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_834 = bc_pe_834_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_835 = bc_pe_835_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_836 = bc_pe_836_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_837 = bc_pe_837_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_838 = bc_pe_838_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_839 = bc_pe_839_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_840 = bc_pe_840_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_841 = bc_pe_841_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_842 = bc_pe_842_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_843 = bc_pe_843_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_844 = bc_pe_844_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_845 = bc_pe_845_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_846 = bc_pe_846_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_847 = bc_pe_847_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_848 = bc_pe_848_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_849 = bc_pe_849_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_850 = bc_pe_850_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_851 = bc_pe_851_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_852 = bc_pe_852_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_853 = bc_pe_853_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_854 = bc_pe_854_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_855 = bc_pe_855_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_856 = bc_pe_856_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_857 = bc_pe_857_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_858 = bc_pe_858_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_859 = bc_pe_859_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_860 = bc_pe_860_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_861 = bc_pe_861_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_862 = bc_pe_862_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_863 = bc_pe_863_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_864 = bc_pe_864_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_865 = bc_pe_865_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_866 = bc_pe_866_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_867 = bc_pe_867_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_868 = bc_pe_868_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_869 = bc_pe_869_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_870 = bc_pe_870_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_871 = bc_pe_871_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_872 = bc_pe_872_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_873 = bc_pe_873_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_874 = bc_pe_874_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_875 = bc_pe_875_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_876 = bc_pe_876_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_877 = bc_pe_877_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_878 = bc_pe_878_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_879 = bc_pe_879_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_880 = bc_pe_880_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_881 = bc_pe_881_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_882 = bc_pe_882_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_883 = bc_pe_883_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_884 = bc_pe_884_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_885 = bc_pe_885_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_886 = bc_pe_886_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_887 = bc_pe_887_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_888 = bc_pe_888_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_889 = bc_pe_889_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_890 = bc_pe_890_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_891 = bc_pe_891_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_892 = bc_pe_892_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_893 = bc_pe_893_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_894 = bc_pe_894_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_895 = bc_pe_895_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_896 = bc_pe_896_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_897 = bc_pe_897_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_898 = bc_pe_898_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_899 = bc_pe_899_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_900 = bc_pe_900_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_901 = bc_pe_901_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_902 = bc_pe_902_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_903 = bc_pe_903_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_904 = bc_pe_904_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_905 = bc_pe_905_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_906 = bc_pe_906_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_907 = bc_pe_907_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_908 = bc_pe_908_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_909 = bc_pe_909_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_910 = bc_pe_910_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_911 = bc_pe_911_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_912 = bc_pe_912_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_913 = bc_pe_913_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_914 = bc_pe_914_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_915 = bc_pe_915_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_916 = bc_pe_916_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_917 = bc_pe_917_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_918 = bc_pe_918_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_919 = bc_pe_919_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_920 = bc_pe_920_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_921 = bc_pe_921_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_922 = bc_pe_922_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_923 = bc_pe_923_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_924 = bc_pe_924_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_925 = bc_pe_925_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_926 = bc_pe_926_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_927 = bc_pe_927_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_928 = bc_pe_928_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_929 = bc_pe_929_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_930 = bc_pe_930_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_931 = bc_pe_931_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_932 = bc_pe_932_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_933 = bc_pe_933_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_934 = bc_pe_934_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_935 = bc_pe_935_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_936 = bc_pe_936_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_937 = bc_pe_937_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_938 = bc_pe_938_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_939 = bc_pe_939_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_940 = bc_pe_940_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_941 = bc_pe_941_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_942 = bc_pe_942_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_943 = bc_pe_943_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_944 = bc_pe_944_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_945 = bc_pe_945_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_946 = bc_pe_946_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_947 = bc_pe_947_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_948 = bc_pe_948_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_949 = bc_pe_949_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_950 = bc_pe_950_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_951 = bc_pe_951_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_952 = bc_pe_952_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_953 = bc_pe_953_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_954 = bc_pe_954_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_955 = bc_pe_955_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_956 = bc_pe_956_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_957 = bc_pe_957_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_958 = bc_pe_958_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_959 = bc_pe_959_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_960 = bc_pe_960_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_961 = bc_pe_961_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_962 = bc_pe_962_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_963 = bc_pe_963_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_964 = bc_pe_964_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_965 = bc_pe_965_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_966 = bc_pe_966_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_967 = bc_pe_967_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_968 = bc_pe_968_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_969 = bc_pe_969_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_970 = bc_pe_970_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_971 = bc_pe_971_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_972 = bc_pe_972_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_973 = bc_pe_973_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_974 = bc_pe_974_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_975 = bc_pe_975_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_976 = bc_pe_976_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_977 = bc_pe_977_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_978 = bc_pe_978_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_979 = bc_pe_979_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_980 = bc_pe_980_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_981 = bc_pe_981_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_982 = bc_pe_982_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_983 = bc_pe_983_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_984 = bc_pe_984_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_985 = bc_pe_985_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_986 = bc_pe_986_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_987 = bc_pe_987_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_988 = bc_pe_988_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_989 = bc_pe_989_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_990 = bc_pe_990_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_991 = bc_pe_991_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_992 = bc_pe_992_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_993 = bc_pe_993_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_994 = bc_pe_994_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_995 = bc_pe_995_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_996 = bc_pe_996_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_997 = bc_pe_997_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_998 = bc_pe_998_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_999 = bc_pe_999_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1000 = bc_pe_1000_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1001 = bc_pe_1001_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1002 = bc_pe_1002_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1003 = bc_pe_1003_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1004 = bc_pe_1004_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1005 = bc_pe_1005_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1006 = bc_pe_1006_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1007 = bc_pe_1007_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1008 = bc_pe_1008_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1009 = bc_pe_1009_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1010 = bc_pe_1010_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1011 = bc_pe_1011_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1012 = bc_pe_1012_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1013 = bc_pe_1013_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1014 = bc_pe_1014_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1015 = bc_pe_1015_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1016 = bc_pe_1016_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1017 = bc_pe_1017_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1018 = bc_pe_1018_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1019 = bc_pe_1019_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1020 = bc_pe_1020_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1021 = bc_pe_1021_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1022 = bc_pe_1022_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1023 = bc_pe_1023_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_clock = clock;
  assign bc_pe_reset = reset;
  assign bc_pe_io_ho_input = io_x_input_0; // @[bc_mmul.scala 22:28 38:42]
  assign bc_pe_io_ve_input = io_w_input_0; // @[bc_mmul.scala 22:28 37:42]
  assign bc_pe_io_input_valid = io_input_valid_0; // @[bc_mmul.scala 22:28 39:42]
  assign bc_pe_io_iormac = io_iormac_0; // @[bc_mmul.scala 22:28 40:42]
  assign bc_pe_1_clock = clock;
  assign bc_pe_1_reset = reset;
  assign bc_pe_1_io_ho_input = bc_pe_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1_io_ve_input = io_w_input_1; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_1_io_input_valid = io_input_valid_1; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_1_io_iormac = io_iormac_1; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_2_clock = clock;
  assign bc_pe_2_reset = reset;
  assign bc_pe_2_io_ho_input = bc_pe_1_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_2_io_ve_input = io_w_input_2; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_2_io_input_valid = io_input_valid_2; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_2_io_iormac = io_iormac_2; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_3_clock = clock;
  assign bc_pe_3_reset = reset;
  assign bc_pe_3_io_ho_input = bc_pe_2_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_3_io_ve_input = io_w_input_3; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_3_io_input_valid = io_input_valid_3; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_3_io_iormac = io_iormac_3; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_4_clock = clock;
  assign bc_pe_4_reset = reset;
  assign bc_pe_4_io_ho_input = bc_pe_3_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_4_io_ve_input = io_w_input_4; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_4_io_input_valid = io_input_valid_4; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_4_io_iormac = io_iormac_4; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_5_clock = clock;
  assign bc_pe_5_reset = reset;
  assign bc_pe_5_io_ho_input = bc_pe_4_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_5_io_ve_input = io_w_input_5; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_5_io_input_valid = io_input_valid_5; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_5_io_iormac = io_iormac_5; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_6_clock = clock;
  assign bc_pe_6_reset = reset;
  assign bc_pe_6_io_ho_input = bc_pe_5_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_6_io_ve_input = io_w_input_6; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_6_io_input_valid = io_input_valid_6; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_6_io_iormac = io_iormac_6; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_7_clock = clock;
  assign bc_pe_7_reset = reset;
  assign bc_pe_7_io_ho_input = bc_pe_6_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_7_io_ve_input = io_w_input_7; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_7_io_input_valid = io_input_valid_7; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_7_io_iormac = io_iormac_7; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_8_clock = clock;
  assign bc_pe_8_reset = reset;
  assign bc_pe_8_io_ho_input = bc_pe_7_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_8_io_ve_input = io_w_input_8; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_8_io_input_valid = io_input_valid_8; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_8_io_iormac = io_iormac_8; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_9_clock = clock;
  assign bc_pe_9_reset = reset;
  assign bc_pe_9_io_ho_input = bc_pe_8_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_9_io_ve_input = io_w_input_9; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_9_io_input_valid = io_input_valid_9; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_9_io_iormac = io_iormac_9; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_10_clock = clock;
  assign bc_pe_10_reset = reset;
  assign bc_pe_10_io_ho_input = bc_pe_9_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_10_io_ve_input = io_w_input_10; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_10_io_input_valid = io_input_valid_10; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_10_io_iormac = io_iormac_10; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_11_clock = clock;
  assign bc_pe_11_reset = reset;
  assign bc_pe_11_io_ho_input = bc_pe_10_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_11_io_ve_input = io_w_input_11; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_11_io_input_valid = io_input_valid_11; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_11_io_iormac = io_iormac_11; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_12_clock = clock;
  assign bc_pe_12_reset = reset;
  assign bc_pe_12_io_ho_input = bc_pe_11_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_12_io_ve_input = io_w_input_12; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_12_io_input_valid = io_input_valid_12; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_12_io_iormac = io_iormac_12; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_13_clock = clock;
  assign bc_pe_13_reset = reset;
  assign bc_pe_13_io_ho_input = bc_pe_12_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_13_io_ve_input = io_w_input_13; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_13_io_input_valid = io_input_valid_13; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_13_io_iormac = io_iormac_13; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_14_clock = clock;
  assign bc_pe_14_reset = reset;
  assign bc_pe_14_io_ho_input = bc_pe_13_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_14_io_ve_input = io_w_input_14; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_14_io_input_valid = io_input_valid_14; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_14_io_iormac = io_iormac_14; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_15_clock = clock;
  assign bc_pe_15_reset = reset;
  assign bc_pe_15_io_ho_input = bc_pe_14_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_15_io_ve_input = io_w_input_15; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_15_io_input_valid = io_input_valid_15; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_15_io_iormac = io_iormac_15; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_16_clock = clock;
  assign bc_pe_16_reset = reset;
  assign bc_pe_16_io_ho_input = bc_pe_15_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_16_io_ve_input = io_w_input_16; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_16_io_input_valid = io_input_valid_16; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_16_io_iormac = io_iormac_16; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_17_clock = clock;
  assign bc_pe_17_reset = reset;
  assign bc_pe_17_io_ho_input = bc_pe_16_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_17_io_ve_input = io_w_input_17; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_17_io_input_valid = io_input_valid_17; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_17_io_iormac = io_iormac_17; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_18_clock = clock;
  assign bc_pe_18_reset = reset;
  assign bc_pe_18_io_ho_input = bc_pe_17_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_18_io_ve_input = io_w_input_18; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_18_io_input_valid = io_input_valid_18; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_18_io_iormac = io_iormac_18; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_19_clock = clock;
  assign bc_pe_19_reset = reset;
  assign bc_pe_19_io_ho_input = bc_pe_18_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_19_io_ve_input = io_w_input_19; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_19_io_input_valid = io_input_valid_19; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_19_io_iormac = io_iormac_19; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_20_clock = clock;
  assign bc_pe_20_reset = reset;
  assign bc_pe_20_io_ho_input = bc_pe_19_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_20_io_ve_input = io_w_input_20; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_20_io_input_valid = io_input_valid_20; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_20_io_iormac = io_iormac_20; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_21_clock = clock;
  assign bc_pe_21_reset = reset;
  assign bc_pe_21_io_ho_input = bc_pe_20_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_21_io_ve_input = io_w_input_21; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_21_io_input_valid = io_input_valid_21; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_21_io_iormac = io_iormac_21; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_22_clock = clock;
  assign bc_pe_22_reset = reset;
  assign bc_pe_22_io_ho_input = bc_pe_21_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_22_io_ve_input = io_w_input_22; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_22_io_input_valid = io_input_valid_22; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_22_io_iormac = io_iormac_22; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_23_clock = clock;
  assign bc_pe_23_reset = reset;
  assign bc_pe_23_io_ho_input = bc_pe_22_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_23_io_ve_input = io_w_input_23; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_23_io_input_valid = io_input_valid_23; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_23_io_iormac = io_iormac_23; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_24_clock = clock;
  assign bc_pe_24_reset = reset;
  assign bc_pe_24_io_ho_input = bc_pe_23_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_24_io_ve_input = io_w_input_24; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_24_io_input_valid = io_input_valid_24; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_24_io_iormac = io_iormac_24; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_25_clock = clock;
  assign bc_pe_25_reset = reset;
  assign bc_pe_25_io_ho_input = bc_pe_24_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_25_io_ve_input = io_w_input_25; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_25_io_input_valid = io_input_valid_25; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_25_io_iormac = io_iormac_25; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_26_clock = clock;
  assign bc_pe_26_reset = reset;
  assign bc_pe_26_io_ho_input = bc_pe_25_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_26_io_ve_input = io_w_input_26; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_26_io_input_valid = io_input_valid_26; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_26_io_iormac = io_iormac_26; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_27_clock = clock;
  assign bc_pe_27_reset = reset;
  assign bc_pe_27_io_ho_input = bc_pe_26_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_27_io_ve_input = io_w_input_27; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_27_io_input_valid = io_input_valid_27; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_27_io_iormac = io_iormac_27; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_28_clock = clock;
  assign bc_pe_28_reset = reset;
  assign bc_pe_28_io_ho_input = bc_pe_27_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_28_io_ve_input = io_w_input_28; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_28_io_input_valid = io_input_valid_28; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_28_io_iormac = io_iormac_28; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_29_clock = clock;
  assign bc_pe_29_reset = reset;
  assign bc_pe_29_io_ho_input = bc_pe_28_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_29_io_ve_input = io_w_input_29; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_29_io_input_valid = io_input_valid_29; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_29_io_iormac = io_iormac_29; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_30_clock = clock;
  assign bc_pe_30_reset = reset;
  assign bc_pe_30_io_ho_input = bc_pe_29_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_30_io_ve_input = io_w_input_30; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_30_io_input_valid = io_input_valid_30; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_30_io_iormac = io_iormac_30; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_31_clock = clock;
  assign bc_pe_31_reset = reset;
  assign bc_pe_31_io_ho_input = bc_pe_30_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_31_io_ve_input = io_w_input_31; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_31_io_input_valid = io_input_valid_31; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_31_io_iormac = io_iormac_31; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_32_clock = clock;
  assign bc_pe_32_reset = reset;
  assign bc_pe_32_io_ho_input = io_x_input_1; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_32_io_ve_input = bc_pe_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_32_io_input_valid = io_input_valid_32; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_32_io_iormac = io_iormac_32; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_33_clock = clock;
  assign bc_pe_33_reset = reset;
  assign bc_pe_33_io_ho_input = bc_pe_32_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_33_io_ve_input = bc_pe_1_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_33_io_input_valid = io_input_valid_33; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_33_io_iormac = io_iormac_33; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_34_clock = clock;
  assign bc_pe_34_reset = reset;
  assign bc_pe_34_io_ho_input = bc_pe_33_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_34_io_ve_input = bc_pe_2_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_34_io_input_valid = io_input_valid_34; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_34_io_iormac = io_iormac_34; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_35_clock = clock;
  assign bc_pe_35_reset = reset;
  assign bc_pe_35_io_ho_input = bc_pe_34_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_35_io_ve_input = bc_pe_3_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_35_io_input_valid = io_input_valid_35; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_35_io_iormac = io_iormac_35; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_36_clock = clock;
  assign bc_pe_36_reset = reset;
  assign bc_pe_36_io_ho_input = bc_pe_35_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_36_io_ve_input = bc_pe_4_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_36_io_input_valid = io_input_valid_36; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_36_io_iormac = io_iormac_36; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_37_clock = clock;
  assign bc_pe_37_reset = reset;
  assign bc_pe_37_io_ho_input = bc_pe_36_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_37_io_ve_input = bc_pe_5_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_37_io_input_valid = io_input_valid_37; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_37_io_iormac = io_iormac_37; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_38_clock = clock;
  assign bc_pe_38_reset = reset;
  assign bc_pe_38_io_ho_input = bc_pe_37_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_38_io_ve_input = bc_pe_6_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_38_io_input_valid = io_input_valid_38; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_38_io_iormac = io_iormac_38; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_39_clock = clock;
  assign bc_pe_39_reset = reset;
  assign bc_pe_39_io_ho_input = bc_pe_38_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_39_io_ve_input = bc_pe_7_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_39_io_input_valid = io_input_valid_39; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_39_io_iormac = io_iormac_39; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_40_clock = clock;
  assign bc_pe_40_reset = reset;
  assign bc_pe_40_io_ho_input = bc_pe_39_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_40_io_ve_input = bc_pe_8_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_40_io_input_valid = io_input_valid_40; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_40_io_iormac = io_iormac_40; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_41_clock = clock;
  assign bc_pe_41_reset = reset;
  assign bc_pe_41_io_ho_input = bc_pe_40_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_41_io_ve_input = bc_pe_9_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_41_io_input_valid = io_input_valid_41; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_41_io_iormac = io_iormac_41; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_42_clock = clock;
  assign bc_pe_42_reset = reset;
  assign bc_pe_42_io_ho_input = bc_pe_41_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_42_io_ve_input = bc_pe_10_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_42_io_input_valid = io_input_valid_42; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_42_io_iormac = io_iormac_42; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_43_clock = clock;
  assign bc_pe_43_reset = reset;
  assign bc_pe_43_io_ho_input = bc_pe_42_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_43_io_ve_input = bc_pe_11_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_43_io_input_valid = io_input_valid_43; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_43_io_iormac = io_iormac_43; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_44_clock = clock;
  assign bc_pe_44_reset = reset;
  assign bc_pe_44_io_ho_input = bc_pe_43_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_44_io_ve_input = bc_pe_12_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_44_io_input_valid = io_input_valid_44; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_44_io_iormac = io_iormac_44; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_45_clock = clock;
  assign bc_pe_45_reset = reset;
  assign bc_pe_45_io_ho_input = bc_pe_44_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_45_io_ve_input = bc_pe_13_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_45_io_input_valid = io_input_valid_45; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_45_io_iormac = io_iormac_45; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_46_clock = clock;
  assign bc_pe_46_reset = reset;
  assign bc_pe_46_io_ho_input = bc_pe_45_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_46_io_ve_input = bc_pe_14_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_46_io_input_valid = io_input_valid_46; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_46_io_iormac = io_iormac_46; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_47_clock = clock;
  assign bc_pe_47_reset = reset;
  assign bc_pe_47_io_ho_input = bc_pe_46_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_47_io_ve_input = bc_pe_15_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_47_io_input_valid = io_input_valid_47; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_47_io_iormac = io_iormac_47; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_48_clock = clock;
  assign bc_pe_48_reset = reset;
  assign bc_pe_48_io_ho_input = bc_pe_47_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_48_io_ve_input = bc_pe_16_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_48_io_input_valid = io_input_valid_48; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_48_io_iormac = io_iormac_48; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_49_clock = clock;
  assign bc_pe_49_reset = reset;
  assign bc_pe_49_io_ho_input = bc_pe_48_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_49_io_ve_input = bc_pe_17_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_49_io_input_valid = io_input_valid_49; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_49_io_iormac = io_iormac_49; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_50_clock = clock;
  assign bc_pe_50_reset = reset;
  assign bc_pe_50_io_ho_input = bc_pe_49_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_50_io_ve_input = bc_pe_18_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_50_io_input_valid = io_input_valid_50; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_50_io_iormac = io_iormac_50; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_51_clock = clock;
  assign bc_pe_51_reset = reset;
  assign bc_pe_51_io_ho_input = bc_pe_50_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_51_io_ve_input = bc_pe_19_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_51_io_input_valid = io_input_valid_51; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_51_io_iormac = io_iormac_51; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_52_clock = clock;
  assign bc_pe_52_reset = reset;
  assign bc_pe_52_io_ho_input = bc_pe_51_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_52_io_ve_input = bc_pe_20_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_52_io_input_valid = io_input_valid_52; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_52_io_iormac = io_iormac_52; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_53_clock = clock;
  assign bc_pe_53_reset = reset;
  assign bc_pe_53_io_ho_input = bc_pe_52_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_53_io_ve_input = bc_pe_21_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_53_io_input_valid = io_input_valid_53; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_53_io_iormac = io_iormac_53; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_54_clock = clock;
  assign bc_pe_54_reset = reset;
  assign bc_pe_54_io_ho_input = bc_pe_53_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_54_io_ve_input = bc_pe_22_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_54_io_input_valid = io_input_valid_54; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_54_io_iormac = io_iormac_54; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_55_clock = clock;
  assign bc_pe_55_reset = reset;
  assign bc_pe_55_io_ho_input = bc_pe_54_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_55_io_ve_input = bc_pe_23_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_55_io_input_valid = io_input_valid_55; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_55_io_iormac = io_iormac_55; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_56_clock = clock;
  assign bc_pe_56_reset = reset;
  assign bc_pe_56_io_ho_input = bc_pe_55_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_56_io_ve_input = bc_pe_24_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_56_io_input_valid = io_input_valid_56; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_56_io_iormac = io_iormac_56; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_57_clock = clock;
  assign bc_pe_57_reset = reset;
  assign bc_pe_57_io_ho_input = bc_pe_56_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_57_io_ve_input = bc_pe_25_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_57_io_input_valid = io_input_valid_57; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_57_io_iormac = io_iormac_57; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_58_clock = clock;
  assign bc_pe_58_reset = reset;
  assign bc_pe_58_io_ho_input = bc_pe_57_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_58_io_ve_input = bc_pe_26_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_58_io_input_valid = io_input_valid_58; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_58_io_iormac = io_iormac_58; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_59_clock = clock;
  assign bc_pe_59_reset = reset;
  assign bc_pe_59_io_ho_input = bc_pe_58_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_59_io_ve_input = bc_pe_27_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_59_io_input_valid = io_input_valid_59; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_59_io_iormac = io_iormac_59; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_60_clock = clock;
  assign bc_pe_60_reset = reset;
  assign bc_pe_60_io_ho_input = bc_pe_59_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_60_io_ve_input = bc_pe_28_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_60_io_input_valid = io_input_valid_60; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_60_io_iormac = io_iormac_60; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_61_clock = clock;
  assign bc_pe_61_reset = reset;
  assign bc_pe_61_io_ho_input = bc_pe_60_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_61_io_ve_input = bc_pe_29_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_61_io_input_valid = io_input_valid_61; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_61_io_iormac = io_iormac_61; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_62_clock = clock;
  assign bc_pe_62_reset = reset;
  assign bc_pe_62_io_ho_input = bc_pe_61_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_62_io_ve_input = bc_pe_30_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_62_io_input_valid = io_input_valid_62; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_62_io_iormac = io_iormac_62; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_63_clock = clock;
  assign bc_pe_63_reset = reset;
  assign bc_pe_63_io_ho_input = bc_pe_62_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_63_io_ve_input = bc_pe_31_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_63_io_input_valid = io_input_valid_63; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_63_io_iormac = io_iormac_63; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_64_clock = clock;
  assign bc_pe_64_reset = reset;
  assign bc_pe_64_io_ho_input = io_x_input_2; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_64_io_ve_input = bc_pe_32_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_64_io_input_valid = io_input_valid_64; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_64_io_iormac = io_iormac_64; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_65_clock = clock;
  assign bc_pe_65_reset = reset;
  assign bc_pe_65_io_ho_input = bc_pe_64_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_65_io_ve_input = bc_pe_33_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_65_io_input_valid = io_input_valid_65; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_65_io_iormac = io_iormac_65; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_66_clock = clock;
  assign bc_pe_66_reset = reset;
  assign bc_pe_66_io_ho_input = bc_pe_65_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_66_io_ve_input = bc_pe_34_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_66_io_input_valid = io_input_valid_66; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_66_io_iormac = io_iormac_66; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_67_clock = clock;
  assign bc_pe_67_reset = reset;
  assign bc_pe_67_io_ho_input = bc_pe_66_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_67_io_ve_input = bc_pe_35_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_67_io_input_valid = io_input_valid_67; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_67_io_iormac = io_iormac_67; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_68_clock = clock;
  assign bc_pe_68_reset = reset;
  assign bc_pe_68_io_ho_input = bc_pe_67_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_68_io_ve_input = bc_pe_36_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_68_io_input_valid = io_input_valid_68; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_68_io_iormac = io_iormac_68; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_69_clock = clock;
  assign bc_pe_69_reset = reset;
  assign bc_pe_69_io_ho_input = bc_pe_68_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_69_io_ve_input = bc_pe_37_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_69_io_input_valid = io_input_valid_69; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_69_io_iormac = io_iormac_69; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_70_clock = clock;
  assign bc_pe_70_reset = reset;
  assign bc_pe_70_io_ho_input = bc_pe_69_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_70_io_ve_input = bc_pe_38_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_70_io_input_valid = io_input_valid_70; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_70_io_iormac = io_iormac_70; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_71_clock = clock;
  assign bc_pe_71_reset = reset;
  assign bc_pe_71_io_ho_input = bc_pe_70_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_71_io_ve_input = bc_pe_39_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_71_io_input_valid = io_input_valid_71; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_71_io_iormac = io_iormac_71; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_72_clock = clock;
  assign bc_pe_72_reset = reset;
  assign bc_pe_72_io_ho_input = bc_pe_71_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_72_io_ve_input = bc_pe_40_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_72_io_input_valid = io_input_valid_72; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_72_io_iormac = io_iormac_72; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_73_clock = clock;
  assign bc_pe_73_reset = reset;
  assign bc_pe_73_io_ho_input = bc_pe_72_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_73_io_ve_input = bc_pe_41_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_73_io_input_valid = io_input_valid_73; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_73_io_iormac = io_iormac_73; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_74_clock = clock;
  assign bc_pe_74_reset = reset;
  assign bc_pe_74_io_ho_input = bc_pe_73_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_74_io_ve_input = bc_pe_42_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_74_io_input_valid = io_input_valid_74; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_74_io_iormac = io_iormac_74; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_75_clock = clock;
  assign bc_pe_75_reset = reset;
  assign bc_pe_75_io_ho_input = bc_pe_74_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_75_io_ve_input = bc_pe_43_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_75_io_input_valid = io_input_valid_75; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_75_io_iormac = io_iormac_75; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_76_clock = clock;
  assign bc_pe_76_reset = reset;
  assign bc_pe_76_io_ho_input = bc_pe_75_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_76_io_ve_input = bc_pe_44_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_76_io_input_valid = io_input_valid_76; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_76_io_iormac = io_iormac_76; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_77_clock = clock;
  assign bc_pe_77_reset = reset;
  assign bc_pe_77_io_ho_input = bc_pe_76_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_77_io_ve_input = bc_pe_45_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_77_io_input_valid = io_input_valid_77; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_77_io_iormac = io_iormac_77; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_78_clock = clock;
  assign bc_pe_78_reset = reset;
  assign bc_pe_78_io_ho_input = bc_pe_77_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_78_io_ve_input = bc_pe_46_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_78_io_input_valid = io_input_valid_78; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_78_io_iormac = io_iormac_78; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_79_clock = clock;
  assign bc_pe_79_reset = reset;
  assign bc_pe_79_io_ho_input = bc_pe_78_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_79_io_ve_input = bc_pe_47_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_79_io_input_valid = io_input_valid_79; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_79_io_iormac = io_iormac_79; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_80_clock = clock;
  assign bc_pe_80_reset = reset;
  assign bc_pe_80_io_ho_input = bc_pe_79_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_80_io_ve_input = bc_pe_48_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_80_io_input_valid = io_input_valid_80; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_80_io_iormac = io_iormac_80; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_81_clock = clock;
  assign bc_pe_81_reset = reset;
  assign bc_pe_81_io_ho_input = bc_pe_80_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_81_io_ve_input = bc_pe_49_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_81_io_input_valid = io_input_valid_81; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_81_io_iormac = io_iormac_81; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_82_clock = clock;
  assign bc_pe_82_reset = reset;
  assign bc_pe_82_io_ho_input = bc_pe_81_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_82_io_ve_input = bc_pe_50_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_82_io_input_valid = io_input_valid_82; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_82_io_iormac = io_iormac_82; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_83_clock = clock;
  assign bc_pe_83_reset = reset;
  assign bc_pe_83_io_ho_input = bc_pe_82_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_83_io_ve_input = bc_pe_51_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_83_io_input_valid = io_input_valid_83; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_83_io_iormac = io_iormac_83; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_84_clock = clock;
  assign bc_pe_84_reset = reset;
  assign bc_pe_84_io_ho_input = bc_pe_83_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_84_io_ve_input = bc_pe_52_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_84_io_input_valid = io_input_valid_84; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_84_io_iormac = io_iormac_84; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_85_clock = clock;
  assign bc_pe_85_reset = reset;
  assign bc_pe_85_io_ho_input = bc_pe_84_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_85_io_ve_input = bc_pe_53_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_85_io_input_valid = io_input_valid_85; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_85_io_iormac = io_iormac_85; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_86_clock = clock;
  assign bc_pe_86_reset = reset;
  assign bc_pe_86_io_ho_input = bc_pe_85_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_86_io_ve_input = bc_pe_54_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_86_io_input_valid = io_input_valid_86; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_86_io_iormac = io_iormac_86; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_87_clock = clock;
  assign bc_pe_87_reset = reset;
  assign bc_pe_87_io_ho_input = bc_pe_86_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_87_io_ve_input = bc_pe_55_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_87_io_input_valid = io_input_valid_87; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_87_io_iormac = io_iormac_87; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_88_clock = clock;
  assign bc_pe_88_reset = reset;
  assign bc_pe_88_io_ho_input = bc_pe_87_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_88_io_ve_input = bc_pe_56_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_88_io_input_valid = io_input_valid_88; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_88_io_iormac = io_iormac_88; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_89_clock = clock;
  assign bc_pe_89_reset = reset;
  assign bc_pe_89_io_ho_input = bc_pe_88_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_89_io_ve_input = bc_pe_57_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_89_io_input_valid = io_input_valid_89; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_89_io_iormac = io_iormac_89; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_90_clock = clock;
  assign bc_pe_90_reset = reset;
  assign bc_pe_90_io_ho_input = bc_pe_89_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_90_io_ve_input = bc_pe_58_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_90_io_input_valid = io_input_valid_90; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_90_io_iormac = io_iormac_90; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_91_clock = clock;
  assign bc_pe_91_reset = reset;
  assign bc_pe_91_io_ho_input = bc_pe_90_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_91_io_ve_input = bc_pe_59_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_91_io_input_valid = io_input_valid_91; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_91_io_iormac = io_iormac_91; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_92_clock = clock;
  assign bc_pe_92_reset = reset;
  assign bc_pe_92_io_ho_input = bc_pe_91_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_92_io_ve_input = bc_pe_60_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_92_io_input_valid = io_input_valid_92; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_92_io_iormac = io_iormac_92; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_93_clock = clock;
  assign bc_pe_93_reset = reset;
  assign bc_pe_93_io_ho_input = bc_pe_92_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_93_io_ve_input = bc_pe_61_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_93_io_input_valid = io_input_valid_93; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_93_io_iormac = io_iormac_93; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_94_clock = clock;
  assign bc_pe_94_reset = reset;
  assign bc_pe_94_io_ho_input = bc_pe_93_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_94_io_ve_input = bc_pe_62_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_94_io_input_valid = io_input_valid_94; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_94_io_iormac = io_iormac_94; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_95_clock = clock;
  assign bc_pe_95_reset = reset;
  assign bc_pe_95_io_ho_input = bc_pe_94_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_95_io_ve_input = bc_pe_63_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_95_io_input_valid = io_input_valid_95; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_95_io_iormac = io_iormac_95; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_96_clock = clock;
  assign bc_pe_96_reset = reset;
  assign bc_pe_96_io_ho_input = io_x_input_3; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_96_io_ve_input = bc_pe_64_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_96_io_input_valid = io_input_valid_96; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_96_io_iormac = io_iormac_96; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_97_clock = clock;
  assign bc_pe_97_reset = reset;
  assign bc_pe_97_io_ho_input = bc_pe_96_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_97_io_ve_input = bc_pe_65_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_97_io_input_valid = io_input_valid_97; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_97_io_iormac = io_iormac_97; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_98_clock = clock;
  assign bc_pe_98_reset = reset;
  assign bc_pe_98_io_ho_input = bc_pe_97_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_98_io_ve_input = bc_pe_66_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_98_io_input_valid = io_input_valid_98; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_98_io_iormac = io_iormac_98; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_99_clock = clock;
  assign bc_pe_99_reset = reset;
  assign bc_pe_99_io_ho_input = bc_pe_98_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_99_io_ve_input = bc_pe_67_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_99_io_input_valid = io_input_valid_99; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_99_io_iormac = io_iormac_99; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_100_clock = clock;
  assign bc_pe_100_reset = reset;
  assign bc_pe_100_io_ho_input = bc_pe_99_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_100_io_ve_input = bc_pe_68_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_100_io_input_valid = io_input_valid_100; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_100_io_iormac = io_iormac_100; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_101_clock = clock;
  assign bc_pe_101_reset = reset;
  assign bc_pe_101_io_ho_input = bc_pe_100_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_101_io_ve_input = bc_pe_69_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_101_io_input_valid = io_input_valid_101; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_101_io_iormac = io_iormac_101; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_102_clock = clock;
  assign bc_pe_102_reset = reset;
  assign bc_pe_102_io_ho_input = bc_pe_101_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_102_io_ve_input = bc_pe_70_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_102_io_input_valid = io_input_valid_102; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_102_io_iormac = io_iormac_102; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_103_clock = clock;
  assign bc_pe_103_reset = reset;
  assign bc_pe_103_io_ho_input = bc_pe_102_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_103_io_ve_input = bc_pe_71_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_103_io_input_valid = io_input_valid_103; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_103_io_iormac = io_iormac_103; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_104_clock = clock;
  assign bc_pe_104_reset = reset;
  assign bc_pe_104_io_ho_input = bc_pe_103_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_104_io_ve_input = bc_pe_72_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_104_io_input_valid = io_input_valid_104; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_104_io_iormac = io_iormac_104; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_105_clock = clock;
  assign bc_pe_105_reset = reset;
  assign bc_pe_105_io_ho_input = bc_pe_104_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_105_io_ve_input = bc_pe_73_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_105_io_input_valid = io_input_valid_105; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_105_io_iormac = io_iormac_105; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_106_clock = clock;
  assign bc_pe_106_reset = reset;
  assign bc_pe_106_io_ho_input = bc_pe_105_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_106_io_ve_input = bc_pe_74_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_106_io_input_valid = io_input_valid_106; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_106_io_iormac = io_iormac_106; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_107_clock = clock;
  assign bc_pe_107_reset = reset;
  assign bc_pe_107_io_ho_input = bc_pe_106_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_107_io_ve_input = bc_pe_75_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_107_io_input_valid = io_input_valid_107; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_107_io_iormac = io_iormac_107; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_108_clock = clock;
  assign bc_pe_108_reset = reset;
  assign bc_pe_108_io_ho_input = bc_pe_107_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_108_io_ve_input = bc_pe_76_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_108_io_input_valid = io_input_valid_108; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_108_io_iormac = io_iormac_108; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_109_clock = clock;
  assign bc_pe_109_reset = reset;
  assign bc_pe_109_io_ho_input = bc_pe_108_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_109_io_ve_input = bc_pe_77_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_109_io_input_valid = io_input_valid_109; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_109_io_iormac = io_iormac_109; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_110_clock = clock;
  assign bc_pe_110_reset = reset;
  assign bc_pe_110_io_ho_input = bc_pe_109_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_110_io_ve_input = bc_pe_78_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_110_io_input_valid = io_input_valid_110; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_110_io_iormac = io_iormac_110; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_111_clock = clock;
  assign bc_pe_111_reset = reset;
  assign bc_pe_111_io_ho_input = bc_pe_110_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_111_io_ve_input = bc_pe_79_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_111_io_input_valid = io_input_valid_111; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_111_io_iormac = io_iormac_111; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_112_clock = clock;
  assign bc_pe_112_reset = reset;
  assign bc_pe_112_io_ho_input = bc_pe_111_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_112_io_ve_input = bc_pe_80_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_112_io_input_valid = io_input_valid_112; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_112_io_iormac = io_iormac_112; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_113_clock = clock;
  assign bc_pe_113_reset = reset;
  assign bc_pe_113_io_ho_input = bc_pe_112_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_113_io_ve_input = bc_pe_81_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_113_io_input_valid = io_input_valid_113; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_113_io_iormac = io_iormac_113; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_114_clock = clock;
  assign bc_pe_114_reset = reset;
  assign bc_pe_114_io_ho_input = bc_pe_113_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_114_io_ve_input = bc_pe_82_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_114_io_input_valid = io_input_valid_114; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_114_io_iormac = io_iormac_114; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_115_clock = clock;
  assign bc_pe_115_reset = reset;
  assign bc_pe_115_io_ho_input = bc_pe_114_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_115_io_ve_input = bc_pe_83_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_115_io_input_valid = io_input_valid_115; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_115_io_iormac = io_iormac_115; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_116_clock = clock;
  assign bc_pe_116_reset = reset;
  assign bc_pe_116_io_ho_input = bc_pe_115_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_116_io_ve_input = bc_pe_84_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_116_io_input_valid = io_input_valid_116; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_116_io_iormac = io_iormac_116; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_117_clock = clock;
  assign bc_pe_117_reset = reset;
  assign bc_pe_117_io_ho_input = bc_pe_116_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_117_io_ve_input = bc_pe_85_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_117_io_input_valid = io_input_valid_117; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_117_io_iormac = io_iormac_117; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_118_clock = clock;
  assign bc_pe_118_reset = reset;
  assign bc_pe_118_io_ho_input = bc_pe_117_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_118_io_ve_input = bc_pe_86_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_118_io_input_valid = io_input_valid_118; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_118_io_iormac = io_iormac_118; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_119_clock = clock;
  assign bc_pe_119_reset = reset;
  assign bc_pe_119_io_ho_input = bc_pe_118_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_119_io_ve_input = bc_pe_87_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_119_io_input_valid = io_input_valid_119; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_119_io_iormac = io_iormac_119; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_120_clock = clock;
  assign bc_pe_120_reset = reset;
  assign bc_pe_120_io_ho_input = bc_pe_119_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_120_io_ve_input = bc_pe_88_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_120_io_input_valid = io_input_valid_120; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_120_io_iormac = io_iormac_120; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_121_clock = clock;
  assign bc_pe_121_reset = reset;
  assign bc_pe_121_io_ho_input = bc_pe_120_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_121_io_ve_input = bc_pe_89_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_121_io_input_valid = io_input_valid_121; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_121_io_iormac = io_iormac_121; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_122_clock = clock;
  assign bc_pe_122_reset = reset;
  assign bc_pe_122_io_ho_input = bc_pe_121_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_122_io_ve_input = bc_pe_90_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_122_io_input_valid = io_input_valid_122; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_122_io_iormac = io_iormac_122; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_123_clock = clock;
  assign bc_pe_123_reset = reset;
  assign bc_pe_123_io_ho_input = bc_pe_122_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_123_io_ve_input = bc_pe_91_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_123_io_input_valid = io_input_valid_123; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_123_io_iormac = io_iormac_123; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_124_clock = clock;
  assign bc_pe_124_reset = reset;
  assign bc_pe_124_io_ho_input = bc_pe_123_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_124_io_ve_input = bc_pe_92_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_124_io_input_valid = io_input_valid_124; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_124_io_iormac = io_iormac_124; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_125_clock = clock;
  assign bc_pe_125_reset = reset;
  assign bc_pe_125_io_ho_input = bc_pe_124_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_125_io_ve_input = bc_pe_93_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_125_io_input_valid = io_input_valid_125; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_125_io_iormac = io_iormac_125; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_126_clock = clock;
  assign bc_pe_126_reset = reset;
  assign bc_pe_126_io_ho_input = bc_pe_125_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_126_io_ve_input = bc_pe_94_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_126_io_input_valid = io_input_valid_126; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_126_io_iormac = io_iormac_126; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_127_clock = clock;
  assign bc_pe_127_reset = reset;
  assign bc_pe_127_io_ho_input = bc_pe_126_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_127_io_ve_input = bc_pe_95_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_127_io_input_valid = io_input_valid_127; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_127_io_iormac = io_iormac_127; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_128_clock = clock;
  assign bc_pe_128_reset = reset;
  assign bc_pe_128_io_ho_input = io_x_input_4; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_128_io_ve_input = bc_pe_96_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_128_io_input_valid = io_input_valid_128; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_128_io_iormac = io_iormac_128; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_129_clock = clock;
  assign bc_pe_129_reset = reset;
  assign bc_pe_129_io_ho_input = bc_pe_128_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_129_io_ve_input = bc_pe_97_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_129_io_input_valid = io_input_valid_129; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_129_io_iormac = io_iormac_129; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_130_clock = clock;
  assign bc_pe_130_reset = reset;
  assign bc_pe_130_io_ho_input = bc_pe_129_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_130_io_ve_input = bc_pe_98_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_130_io_input_valid = io_input_valid_130; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_130_io_iormac = io_iormac_130; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_131_clock = clock;
  assign bc_pe_131_reset = reset;
  assign bc_pe_131_io_ho_input = bc_pe_130_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_131_io_ve_input = bc_pe_99_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_131_io_input_valid = io_input_valid_131; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_131_io_iormac = io_iormac_131; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_132_clock = clock;
  assign bc_pe_132_reset = reset;
  assign bc_pe_132_io_ho_input = bc_pe_131_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_132_io_ve_input = bc_pe_100_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_132_io_input_valid = io_input_valid_132; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_132_io_iormac = io_iormac_132; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_133_clock = clock;
  assign bc_pe_133_reset = reset;
  assign bc_pe_133_io_ho_input = bc_pe_132_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_133_io_ve_input = bc_pe_101_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_133_io_input_valid = io_input_valid_133; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_133_io_iormac = io_iormac_133; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_134_clock = clock;
  assign bc_pe_134_reset = reset;
  assign bc_pe_134_io_ho_input = bc_pe_133_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_134_io_ve_input = bc_pe_102_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_134_io_input_valid = io_input_valid_134; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_134_io_iormac = io_iormac_134; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_135_clock = clock;
  assign bc_pe_135_reset = reset;
  assign bc_pe_135_io_ho_input = bc_pe_134_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_135_io_ve_input = bc_pe_103_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_135_io_input_valid = io_input_valid_135; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_135_io_iormac = io_iormac_135; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_136_clock = clock;
  assign bc_pe_136_reset = reset;
  assign bc_pe_136_io_ho_input = bc_pe_135_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_136_io_ve_input = bc_pe_104_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_136_io_input_valid = io_input_valid_136; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_136_io_iormac = io_iormac_136; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_137_clock = clock;
  assign bc_pe_137_reset = reset;
  assign bc_pe_137_io_ho_input = bc_pe_136_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_137_io_ve_input = bc_pe_105_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_137_io_input_valid = io_input_valid_137; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_137_io_iormac = io_iormac_137; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_138_clock = clock;
  assign bc_pe_138_reset = reset;
  assign bc_pe_138_io_ho_input = bc_pe_137_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_138_io_ve_input = bc_pe_106_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_138_io_input_valid = io_input_valid_138; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_138_io_iormac = io_iormac_138; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_139_clock = clock;
  assign bc_pe_139_reset = reset;
  assign bc_pe_139_io_ho_input = bc_pe_138_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_139_io_ve_input = bc_pe_107_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_139_io_input_valid = io_input_valid_139; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_139_io_iormac = io_iormac_139; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_140_clock = clock;
  assign bc_pe_140_reset = reset;
  assign bc_pe_140_io_ho_input = bc_pe_139_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_140_io_ve_input = bc_pe_108_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_140_io_input_valid = io_input_valid_140; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_140_io_iormac = io_iormac_140; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_141_clock = clock;
  assign bc_pe_141_reset = reset;
  assign bc_pe_141_io_ho_input = bc_pe_140_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_141_io_ve_input = bc_pe_109_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_141_io_input_valid = io_input_valid_141; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_141_io_iormac = io_iormac_141; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_142_clock = clock;
  assign bc_pe_142_reset = reset;
  assign bc_pe_142_io_ho_input = bc_pe_141_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_142_io_ve_input = bc_pe_110_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_142_io_input_valid = io_input_valid_142; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_142_io_iormac = io_iormac_142; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_143_clock = clock;
  assign bc_pe_143_reset = reset;
  assign bc_pe_143_io_ho_input = bc_pe_142_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_143_io_ve_input = bc_pe_111_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_143_io_input_valid = io_input_valid_143; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_143_io_iormac = io_iormac_143; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_144_clock = clock;
  assign bc_pe_144_reset = reset;
  assign bc_pe_144_io_ho_input = bc_pe_143_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_144_io_ve_input = bc_pe_112_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_144_io_input_valid = io_input_valid_144; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_144_io_iormac = io_iormac_144; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_145_clock = clock;
  assign bc_pe_145_reset = reset;
  assign bc_pe_145_io_ho_input = bc_pe_144_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_145_io_ve_input = bc_pe_113_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_145_io_input_valid = io_input_valid_145; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_145_io_iormac = io_iormac_145; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_146_clock = clock;
  assign bc_pe_146_reset = reset;
  assign bc_pe_146_io_ho_input = bc_pe_145_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_146_io_ve_input = bc_pe_114_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_146_io_input_valid = io_input_valid_146; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_146_io_iormac = io_iormac_146; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_147_clock = clock;
  assign bc_pe_147_reset = reset;
  assign bc_pe_147_io_ho_input = bc_pe_146_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_147_io_ve_input = bc_pe_115_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_147_io_input_valid = io_input_valid_147; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_147_io_iormac = io_iormac_147; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_148_clock = clock;
  assign bc_pe_148_reset = reset;
  assign bc_pe_148_io_ho_input = bc_pe_147_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_148_io_ve_input = bc_pe_116_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_148_io_input_valid = io_input_valid_148; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_148_io_iormac = io_iormac_148; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_149_clock = clock;
  assign bc_pe_149_reset = reset;
  assign bc_pe_149_io_ho_input = bc_pe_148_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_149_io_ve_input = bc_pe_117_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_149_io_input_valid = io_input_valid_149; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_149_io_iormac = io_iormac_149; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_150_clock = clock;
  assign bc_pe_150_reset = reset;
  assign bc_pe_150_io_ho_input = bc_pe_149_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_150_io_ve_input = bc_pe_118_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_150_io_input_valid = io_input_valid_150; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_150_io_iormac = io_iormac_150; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_151_clock = clock;
  assign bc_pe_151_reset = reset;
  assign bc_pe_151_io_ho_input = bc_pe_150_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_151_io_ve_input = bc_pe_119_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_151_io_input_valid = io_input_valid_151; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_151_io_iormac = io_iormac_151; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_152_clock = clock;
  assign bc_pe_152_reset = reset;
  assign bc_pe_152_io_ho_input = bc_pe_151_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_152_io_ve_input = bc_pe_120_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_152_io_input_valid = io_input_valid_152; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_152_io_iormac = io_iormac_152; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_153_clock = clock;
  assign bc_pe_153_reset = reset;
  assign bc_pe_153_io_ho_input = bc_pe_152_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_153_io_ve_input = bc_pe_121_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_153_io_input_valid = io_input_valid_153; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_153_io_iormac = io_iormac_153; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_154_clock = clock;
  assign bc_pe_154_reset = reset;
  assign bc_pe_154_io_ho_input = bc_pe_153_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_154_io_ve_input = bc_pe_122_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_154_io_input_valid = io_input_valid_154; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_154_io_iormac = io_iormac_154; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_155_clock = clock;
  assign bc_pe_155_reset = reset;
  assign bc_pe_155_io_ho_input = bc_pe_154_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_155_io_ve_input = bc_pe_123_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_155_io_input_valid = io_input_valid_155; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_155_io_iormac = io_iormac_155; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_156_clock = clock;
  assign bc_pe_156_reset = reset;
  assign bc_pe_156_io_ho_input = bc_pe_155_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_156_io_ve_input = bc_pe_124_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_156_io_input_valid = io_input_valid_156; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_156_io_iormac = io_iormac_156; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_157_clock = clock;
  assign bc_pe_157_reset = reset;
  assign bc_pe_157_io_ho_input = bc_pe_156_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_157_io_ve_input = bc_pe_125_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_157_io_input_valid = io_input_valid_157; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_157_io_iormac = io_iormac_157; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_158_clock = clock;
  assign bc_pe_158_reset = reset;
  assign bc_pe_158_io_ho_input = bc_pe_157_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_158_io_ve_input = bc_pe_126_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_158_io_input_valid = io_input_valid_158; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_158_io_iormac = io_iormac_158; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_159_clock = clock;
  assign bc_pe_159_reset = reset;
  assign bc_pe_159_io_ho_input = bc_pe_158_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_159_io_ve_input = bc_pe_127_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_159_io_input_valid = io_input_valid_159; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_159_io_iormac = io_iormac_159; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_160_clock = clock;
  assign bc_pe_160_reset = reset;
  assign bc_pe_160_io_ho_input = io_x_input_5; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_160_io_ve_input = bc_pe_128_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_160_io_input_valid = io_input_valid_160; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_160_io_iormac = io_iormac_160; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_161_clock = clock;
  assign bc_pe_161_reset = reset;
  assign bc_pe_161_io_ho_input = bc_pe_160_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_161_io_ve_input = bc_pe_129_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_161_io_input_valid = io_input_valid_161; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_161_io_iormac = io_iormac_161; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_162_clock = clock;
  assign bc_pe_162_reset = reset;
  assign bc_pe_162_io_ho_input = bc_pe_161_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_162_io_ve_input = bc_pe_130_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_162_io_input_valid = io_input_valid_162; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_162_io_iormac = io_iormac_162; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_163_clock = clock;
  assign bc_pe_163_reset = reset;
  assign bc_pe_163_io_ho_input = bc_pe_162_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_163_io_ve_input = bc_pe_131_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_163_io_input_valid = io_input_valid_163; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_163_io_iormac = io_iormac_163; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_164_clock = clock;
  assign bc_pe_164_reset = reset;
  assign bc_pe_164_io_ho_input = bc_pe_163_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_164_io_ve_input = bc_pe_132_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_164_io_input_valid = io_input_valid_164; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_164_io_iormac = io_iormac_164; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_165_clock = clock;
  assign bc_pe_165_reset = reset;
  assign bc_pe_165_io_ho_input = bc_pe_164_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_165_io_ve_input = bc_pe_133_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_165_io_input_valid = io_input_valid_165; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_165_io_iormac = io_iormac_165; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_166_clock = clock;
  assign bc_pe_166_reset = reset;
  assign bc_pe_166_io_ho_input = bc_pe_165_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_166_io_ve_input = bc_pe_134_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_166_io_input_valid = io_input_valid_166; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_166_io_iormac = io_iormac_166; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_167_clock = clock;
  assign bc_pe_167_reset = reset;
  assign bc_pe_167_io_ho_input = bc_pe_166_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_167_io_ve_input = bc_pe_135_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_167_io_input_valid = io_input_valid_167; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_167_io_iormac = io_iormac_167; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_168_clock = clock;
  assign bc_pe_168_reset = reset;
  assign bc_pe_168_io_ho_input = bc_pe_167_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_168_io_ve_input = bc_pe_136_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_168_io_input_valid = io_input_valid_168; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_168_io_iormac = io_iormac_168; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_169_clock = clock;
  assign bc_pe_169_reset = reset;
  assign bc_pe_169_io_ho_input = bc_pe_168_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_169_io_ve_input = bc_pe_137_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_169_io_input_valid = io_input_valid_169; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_169_io_iormac = io_iormac_169; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_170_clock = clock;
  assign bc_pe_170_reset = reset;
  assign bc_pe_170_io_ho_input = bc_pe_169_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_170_io_ve_input = bc_pe_138_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_170_io_input_valid = io_input_valid_170; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_170_io_iormac = io_iormac_170; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_171_clock = clock;
  assign bc_pe_171_reset = reset;
  assign bc_pe_171_io_ho_input = bc_pe_170_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_171_io_ve_input = bc_pe_139_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_171_io_input_valid = io_input_valid_171; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_171_io_iormac = io_iormac_171; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_172_clock = clock;
  assign bc_pe_172_reset = reset;
  assign bc_pe_172_io_ho_input = bc_pe_171_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_172_io_ve_input = bc_pe_140_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_172_io_input_valid = io_input_valid_172; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_172_io_iormac = io_iormac_172; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_173_clock = clock;
  assign bc_pe_173_reset = reset;
  assign bc_pe_173_io_ho_input = bc_pe_172_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_173_io_ve_input = bc_pe_141_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_173_io_input_valid = io_input_valid_173; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_173_io_iormac = io_iormac_173; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_174_clock = clock;
  assign bc_pe_174_reset = reset;
  assign bc_pe_174_io_ho_input = bc_pe_173_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_174_io_ve_input = bc_pe_142_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_174_io_input_valid = io_input_valid_174; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_174_io_iormac = io_iormac_174; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_175_clock = clock;
  assign bc_pe_175_reset = reset;
  assign bc_pe_175_io_ho_input = bc_pe_174_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_175_io_ve_input = bc_pe_143_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_175_io_input_valid = io_input_valid_175; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_175_io_iormac = io_iormac_175; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_176_clock = clock;
  assign bc_pe_176_reset = reset;
  assign bc_pe_176_io_ho_input = bc_pe_175_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_176_io_ve_input = bc_pe_144_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_176_io_input_valid = io_input_valid_176; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_176_io_iormac = io_iormac_176; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_177_clock = clock;
  assign bc_pe_177_reset = reset;
  assign bc_pe_177_io_ho_input = bc_pe_176_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_177_io_ve_input = bc_pe_145_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_177_io_input_valid = io_input_valid_177; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_177_io_iormac = io_iormac_177; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_178_clock = clock;
  assign bc_pe_178_reset = reset;
  assign bc_pe_178_io_ho_input = bc_pe_177_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_178_io_ve_input = bc_pe_146_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_178_io_input_valid = io_input_valid_178; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_178_io_iormac = io_iormac_178; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_179_clock = clock;
  assign bc_pe_179_reset = reset;
  assign bc_pe_179_io_ho_input = bc_pe_178_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_179_io_ve_input = bc_pe_147_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_179_io_input_valid = io_input_valid_179; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_179_io_iormac = io_iormac_179; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_180_clock = clock;
  assign bc_pe_180_reset = reset;
  assign bc_pe_180_io_ho_input = bc_pe_179_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_180_io_ve_input = bc_pe_148_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_180_io_input_valid = io_input_valid_180; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_180_io_iormac = io_iormac_180; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_181_clock = clock;
  assign bc_pe_181_reset = reset;
  assign bc_pe_181_io_ho_input = bc_pe_180_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_181_io_ve_input = bc_pe_149_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_181_io_input_valid = io_input_valid_181; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_181_io_iormac = io_iormac_181; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_182_clock = clock;
  assign bc_pe_182_reset = reset;
  assign bc_pe_182_io_ho_input = bc_pe_181_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_182_io_ve_input = bc_pe_150_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_182_io_input_valid = io_input_valid_182; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_182_io_iormac = io_iormac_182; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_183_clock = clock;
  assign bc_pe_183_reset = reset;
  assign bc_pe_183_io_ho_input = bc_pe_182_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_183_io_ve_input = bc_pe_151_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_183_io_input_valid = io_input_valid_183; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_183_io_iormac = io_iormac_183; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_184_clock = clock;
  assign bc_pe_184_reset = reset;
  assign bc_pe_184_io_ho_input = bc_pe_183_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_184_io_ve_input = bc_pe_152_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_184_io_input_valid = io_input_valid_184; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_184_io_iormac = io_iormac_184; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_185_clock = clock;
  assign bc_pe_185_reset = reset;
  assign bc_pe_185_io_ho_input = bc_pe_184_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_185_io_ve_input = bc_pe_153_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_185_io_input_valid = io_input_valid_185; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_185_io_iormac = io_iormac_185; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_186_clock = clock;
  assign bc_pe_186_reset = reset;
  assign bc_pe_186_io_ho_input = bc_pe_185_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_186_io_ve_input = bc_pe_154_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_186_io_input_valid = io_input_valid_186; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_186_io_iormac = io_iormac_186; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_187_clock = clock;
  assign bc_pe_187_reset = reset;
  assign bc_pe_187_io_ho_input = bc_pe_186_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_187_io_ve_input = bc_pe_155_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_187_io_input_valid = io_input_valid_187; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_187_io_iormac = io_iormac_187; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_188_clock = clock;
  assign bc_pe_188_reset = reset;
  assign bc_pe_188_io_ho_input = bc_pe_187_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_188_io_ve_input = bc_pe_156_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_188_io_input_valid = io_input_valid_188; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_188_io_iormac = io_iormac_188; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_189_clock = clock;
  assign bc_pe_189_reset = reset;
  assign bc_pe_189_io_ho_input = bc_pe_188_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_189_io_ve_input = bc_pe_157_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_189_io_input_valid = io_input_valid_189; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_189_io_iormac = io_iormac_189; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_190_clock = clock;
  assign bc_pe_190_reset = reset;
  assign bc_pe_190_io_ho_input = bc_pe_189_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_190_io_ve_input = bc_pe_158_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_190_io_input_valid = io_input_valid_190; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_190_io_iormac = io_iormac_190; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_191_clock = clock;
  assign bc_pe_191_reset = reset;
  assign bc_pe_191_io_ho_input = bc_pe_190_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_191_io_ve_input = bc_pe_159_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_191_io_input_valid = io_input_valid_191; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_191_io_iormac = io_iormac_191; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_192_clock = clock;
  assign bc_pe_192_reset = reset;
  assign bc_pe_192_io_ho_input = io_x_input_6; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_192_io_ve_input = bc_pe_160_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_192_io_input_valid = io_input_valid_192; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_192_io_iormac = io_iormac_192; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_193_clock = clock;
  assign bc_pe_193_reset = reset;
  assign bc_pe_193_io_ho_input = bc_pe_192_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_193_io_ve_input = bc_pe_161_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_193_io_input_valid = io_input_valid_193; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_193_io_iormac = io_iormac_193; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_194_clock = clock;
  assign bc_pe_194_reset = reset;
  assign bc_pe_194_io_ho_input = bc_pe_193_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_194_io_ve_input = bc_pe_162_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_194_io_input_valid = io_input_valid_194; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_194_io_iormac = io_iormac_194; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_195_clock = clock;
  assign bc_pe_195_reset = reset;
  assign bc_pe_195_io_ho_input = bc_pe_194_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_195_io_ve_input = bc_pe_163_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_195_io_input_valid = io_input_valid_195; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_195_io_iormac = io_iormac_195; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_196_clock = clock;
  assign bc_pe_196_reset = reset;
  assign bc_pe_196_io_ho_input = bc_pe_195_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_196_io_ve_input = bc_pe_164_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_196_io_input_valid = io_input_valid_196; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_196_io_iormac = io_iormac_196; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_197_clock = clock;
  assign bc_pe_197_reset = reset;
  assign bc_pe_197_io_ho_input = bc_pe_196_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_197_io_ve_input = bc_pe_165_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_197_io_input_valid = io_input_valid_197; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_197_io_iormac = io_iormac_197; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_198_clock = clock;
  assign bc_pe_198_reset = reset;
  assign bc_pe_198_io_ho_input = bc_pe_197_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_198_io_ve_input = bc_pe_166_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_198_io_input_valid = io_input_valid_198; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_198_io_iormac = io_iormac_198; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_199_clock = clock;
  assign bc_pe_199_reset = reset;
  assign bc_pe_199_io_ho_input = bc_pe_198_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_199_io_ve_input = bc_pe_167_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_199_io_input_valid = io_input_valid_199; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_199_io_iormac = io_iormac_199; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_200_clock = clock;
  assign bc_pe_200_reset = reset;
  assign bc_pe_200_io_ho_input = bc_pe_199_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_200_io_ve_input = bc_pe_168_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_200_io_input_valid = io_input_valid_200; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_200_io_iormac = io_iormac_200; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_201_clock = clock;
  assign bc_pe_201_reset = reset;
  assign bc_pe_201_io_ho_input = bc_pe_200_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_201_io_ve_input = bc_pe_169_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_201_io_input_valid = io_input_valid_201; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_201_io_iormac = io_iormac_201; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_202_clock = clock;
  assign bc_pe_202_reset = reset;
  assign bc_pe_202_io_ho_input = bc_pe_201_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_202_io_ve_input = bc_pe_170_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_202_io_input_valid = io_input_valid_202; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_202_io_iormac = io_iormac_202; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_203_clock = clock;
  assign bc_pe_203_reset = reset;
  assign bc_pe_203_io_ho_input = bc_pe_202_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_203_io_ve_input = bc_pe_171_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_203_io_input_valid = io_input_valid_203; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_203_io_iormac = io_iormac_203; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_204_clock = clock;
  assign bc_pe_204_reset = reset;
  assign bc_pe_204_io_ho_input = bc_pe_203_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_204_io_ve_input = bc_pe_172_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_204_io_input_valid = io_input_valid_204; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_204_io_iormac = io_iormac_204; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_205_clock = clock;
  assign bc_pe_205_reset = reset;
  assign bc_pe_205_io_ho_input = bc_pe_204_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_205_io_ve_input = bc_pe_173_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_205_io_input_valid = io_input_valid_205; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_205_io_iormac = io_iormac_205; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_206_clock = clock;
  assign bc_pe_206_reset = reset;
  assign bc_pe_206_io_ho_input = bc_pe_205_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_206_io_ve_input = bc_pe_174_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_206_io_input_valid = io_input_valid_206; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_206_io_iormac = io_iormac_206; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_207_clock = clock;
  assign bc_pe_207_reset = reset;
  assign bc_pe_207_io_ho_input = bc_pe_206_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_207_io_ve_input = bc_pe_175_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_207_io_input_valid = io_input_valid_207; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_207_io_iormac = io_iormac_207; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_208_clock = clock;
  assign bc_pe_208_reset = reset;
  assign bc_pe_208_io_ho_input = bc_pe_207_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_208_io_ve_input = bc_pe_176_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_208_io_input_valid = io_input_valid_208; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_208_io_iormac = io_iormac_208; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_209_clock = clock;
  assign bc_pe_209_reset = reset;
  assign bc_pe_209_io_ho_input = bc_pe_208_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_209_io_ve_input = bc_pe_177_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_209_io_input_valid = io_input_valid_209; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_209_io_iormac = io_iormac_209; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_210_clock = clock;
  assign bc_pe_210_reset = reset;
  assign bc_pe_210_io_ho_input = bc_pe_209_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_210_io_ve_input = bc_pe_178_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_210_io_input_valid = io_input_valid_210; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_210_io_iormac = io_iormac_210; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_211_clock = clock;
  assign bc_pe_211_reset = reset;
  assign bc_pe_211_io_ho_input = bc_pe_210_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_211_io_ve_input = bc_pe_179_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_211_io_input_valid = io_input_valid_211; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_211_io_iormac = io_iormac_211; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_212_clock = clock;
  assign bc_pe_212_reset = reset;
  assign bc_pe_212_io_ho_input = bc_pe_211_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_212_io_ve_input = bc_pe_180_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_212_io_input_valid = io_input_valid_212; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_212_io_iormac = io_iormac_212; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_213_clock = clock;
  assign bc_pe_213_reset = reset;
  assign bc_pe_213_io_ho_input = bc_pe_212_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_213_io_ve_input = bc_pe_181_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_213_io_input_valid = io_input_valid_213; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_213_io_iormac = io_iormac_213; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_214_clock = clock;
  assign bc_pe_214_reset = reset;
  assign bc_pe_214_io_ho_input = bc_pe_213_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_214_io_ve_input = bc_pe_182_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_214_io_input_valid = io_input_valid_214; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_214_io_iormac = io_iormac_214; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_215_clock = clock;
  assign bc_pe_215_reset = reset;
  assign bc_pe_215_io_ho_input = bc_pe_214_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_215_io_ve_input = bc_pe_183_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_215_io_input_valid = io_input_valid_215; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_215_io_iormac = io_iormac_215; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_216_clock = clock;
  assign bc_pe_216_reset = reset;
  assign bc_pe_216_io_ho_input = bc_pe_215_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_216_io_ve_input = bc_pe_184_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_216_io_input_valid = io_input_valid_216; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_216_io_iormac = io_iormac_216; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_217_clock = clock;
  assign bc_pe_217_reset = reset;
  assign bc_pe_217_io_ho_input = bc_pe_216_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_217_io_ve_input = bc_pe_185_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_217_io_input_valid = io_input_valid_217; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_217_io_iormac = io_iormac_217; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_218_clock = clock;
  assign bc_pe_218_reset = reset;
  assign bc_pe_218_io_ho_input = bc_pe_217_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_218_io_ve_input = bc_pe_186_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_218_io_input_valid = io_input_valid_218; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_218_io_iormac = io_iormac_218; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_219_clock = clock;
  assign bc_pe_219_reset = reset;
  assign bc_pe_219_io_ho_input = bc_pe_218_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_219_io_ve_input = bc_pe_187_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_219_io_input_valid = io_input_valid_219; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_219_io_iormac = io_iormac_219; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_220_clock = clock;
  assign bc_pe_220_reset = reset;
  assign bc_pe_220_io_ho_input = bc_pe_219_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_220_io_ve_input = bc_pe_188_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_220_io_input_valid = io_input_valid_220; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_220_io_iormac = io_iormac_220; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_221_clock = clock;
  assign bc_pe_221_reset = reset;
  assign bc_pe_221_io_ho_input = bc_pe_220_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_221_io_ve_input = bc_pe_189_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_221_io_input_valid = io_input_valid_221; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_221_io_iormac = io_iormac_221; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_222_clock = clock;
  assign bc_pe_222_reset = reset;
  assign bc_pe_222_io_ho_input = bc_pe_221_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_222_io_ve_input = bc_pe_190_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_222_io_input_valid = io_input_valid_222; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_222_io_iormac = io_iormac_222; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_223_clock = clock;
  assign bc_pe_223_reset = reset;
  assign bc_pe_223_io_ho_input = bc_pe_222_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_223_io_ve_input = bc_pe_191_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_223_io_input_valid = io_input_valid_223; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_223_io_iormac = io_iormac_223; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_224_clock = clock;
  assign bc_pe_224_reset = reset;
  assign bc_pe_224_io_ho_input = io_x_input_7; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_224_io_ve_input = bc_pe_192_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_224_io_input_valid = io_input_valid_224; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_224_io_iormac = io_iormac_224; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_225_clock = clock;
  assign bc_pe_225_reset = reset;
  assign bc_pe_225_io_ho_input = bc_pe_224_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_225_io_ve_input = bc_pe_193_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_225_io_input_valid = io_input_valid_225; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_225_io_iormac = io_iormac_225; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_226_clock = clock;
  assign bc_pe_226_reset = reset;
  assign bc_pe_226_io_ho_input = bc_pe_225_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_226_io_ve_input = bc_pe_194_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_226_io_input_valid = io_input_valid_226; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_226_io_iormac = io_iormac_226; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_227_clock = clock;
  assign bc_pe_227_reset = reset;
  assign bc_pe_227_io_ho_input = bc_pe_226_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_227_io_ve_input = bc_pe_195_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_227_io_input_valid = io_input_valid_227; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_227_io_iormac = io_iormac_227; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_228_clock = clock;
  assign bc_pe_228_reset = reset;
  assign bc_pe_228_io_ho_input = bc_pe_227_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_228_io_ve_input = bc_pe_196_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_228_io_input_valid = io_input_valid_228; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_228_io_iormac = io_iormac_228; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_229_clock = clock;
  assign bc_pe_229_reset = reset;
  assign bc_pe_229_io_ho_input = bc_pe_228_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_229_io_ve_input = bc_pe_197_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_229_io_input_valid = io_input_valid_229; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_229_io_iormac = io_iormac_229; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_230_clock = clock;
  assign bc_pe_230_reset = reset;
  assign bc_pe_230_io_ho_input = bc_pe_229_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_230_io_ve_input = bc_pe_198_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_230_io_input_valid = io_input_valid_230; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_230_io_iormac = io_iormac_230; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_231_clock = clock;
  assign bc_pe_231_reset = reset;
  assign bc_pe_231_io_ho_input = bc_pe_230_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_231_io_ve_input = bc_pe_199_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_231_io_input_valid = io_input_valid_231; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_231_io_iormac = io_iormac_231; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_232_clock = clock;
  assign bc_pe_232_reset = reset;
  assign bc_pe_232_io_ho_input = bc_pe_231_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_232_io_ve_input = bc_pe_200_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_232_io_input_valid = io_input_valid_232; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_232_io_iormac = io_iormac_232; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_233_clock = clock;
  assign bc_pe_233_reset = reset;
  assign bc_pe_233_io_ho_input = bc_pe_232_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_233_io_ve_input = bc_pe_201_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_233_io_input_valid = io_input_valid_233; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_233_io_iormac = io_iormac_233; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_234_clock = clock;
  assign bc_pe_234_reset = reset;
  assign bc_pe_234_io_ho_input = bc_pe_233_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_234_io_ve_input = bc_pe_202_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_234_io_input_valid = io_input_valid_234; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_234_io_iormac = io_iormac_234; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_235_clock = clock;
  assign bc_pe_235_reset = reset;
  assign bc_pe_235_io_ho_input = bc_pe_234_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_235_io_ve_input = bc_pe_203_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_235_io_input_valid = io_input_valid_235; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_235_io_iormac = io_iormac_235; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_236_clock = clock;
  assign bc_pe_236_reset = reset;
  assign bc_pe_236_io_ho_input = bc_pe_235_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_236_io_ve_input = bc_pe_204_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_236_io_input_valid = io_input_valid_236; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_236_io_iormac = io_iormac_236; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_237_clock = clock;
  assign bc_pe_237_reset = reset;
  assign bc_pe_237_io_ho_input = bc_pe_236_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_237_io_ve_input = bc_pe_205_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_237_io_input_valid = io_input_valid_237; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_237_io_iormac = io_iormac_237; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_238_clock = clock;
  assign bc_pe_238_reset = reset;
  assign bc_pe_238_io_ho_input = bc_pe_237_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_238_io_ve_input = bc_pe_206_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_238_io_input_valid = io_input_valid_238; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_238_io_iormac = io_iormac_238; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_239_clock = clock;
  assign bc_pe_239_reset = reset;
  assign bc_pe_239_io_ho_input = bc_pe_238_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_239_io_ve_input = bc_pe_207_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_239_io_input_valid = io_input_valid_239; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_239_io_iormac = io_iormac_239; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_240_clock = clock;
  assign bc_pe_240_reset = reset;
  assign bc_pe_240_io_ho_input = bc_pe_239_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_240_io_ve_input = bc_pe_208_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_240_io_input_valid = io_input_valid_240; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_240_io_iormac = io_iormac_240; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_241_clock = clock;
  assign bc_pe_241_reset = reset;
  assign bc_pe_241_io_ho_input = bc_pe_240_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_241_io_ve_input = bc_pe_209_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_241_io_input_valid = io_input_valid_241; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_241_io_iormac = io_iormac_241; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_242_clock = clock;
  assign bc_pe_242_reset = reset;
  assign bc_pe_242_io_ho_input = bc_pe_241_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_242_io_ve_input = bc_pe_210_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_242_io_input_valid = io_input_valid_242; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_242_io_iormac = io_iormac_242; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_243_clock = clock;
  assign bc_pe_243_reset = reset;
  assign bc_pe_243_io_ho_input = bc_pe_242_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_243_io_ve_input = bc_pe_211_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_243_io_input_valid = io_input_valid_243; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_243_io_iormac = io_iormac_243; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_244_clock = clock;
  assign bc_pe_244_reset = reset;
  assign bc_pe_244_io_ho_input = bc_pe_243_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_244_io_ve_input = bc_pe_212_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_244_io_input_valid = io_input_valid_244; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_244_io_iormac = io_iormac_244; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_245_clock = clock;
  assign bc_pe_245_reset = reset;
  assign bc_pe_245_io_ho_input = bc_pe_244_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_245_io_ve_input = bc_pe_213_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_245_io_input_valid = io_input_valid_245; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_245_io_iormac = io_iormac_245; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_246_clock = clock;
  assign bc_pe_246_reset = reset;
  assign bc_pe_246_io_ho_input = bc_pe_245_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_246_io_ve_input = bc_pe_214_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_246_io_input_valid = io_input_valid_246; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_246_io_iormac = io_iormac_246; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_247_clock = clock;
  assign bc_pe_247_reset = reset;
  assign bc_pe_247_io_ho_input = bc_pe_246_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_247_io_ve_input = bc_pe_215_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_247_io_input_valid = io_input_valid_247; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_247_io_iormac = io_iormac_247; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_248_clock = clock;
  assign bc_pe_248_reset = reset;
  assign bc_pe_248_io_ho_input = bc_pe_247_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_248_io_ve_input = bc_pe_216_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_248_io_input_valid = io_input_valid_248; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_248_io_iormac = io_iormac_248; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_249_clock = clock;
  assign bc_pe_249_reset = reset;
  assign bc_pe_249_io_ho_input = bc_pe_248_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_249_io_ve_input = bc_pe_217_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_249_io_input_valid = io_input_valid_249; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_249_io_iormac = io_iormac_249; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_250_clock = clock;
  assign bc_pe_250_reset = reset;
  assign bc_pe_250_io_ho_input = bc_pe_249_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_250_io_ve_input = bc_pe_218_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_250_io_input_valid = io_input_valid_250; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_250_io_iormac = io_iormac_250; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_251_clock = clock;
  assign bc_pe_251_reset = reset;
  assign bc_pe_251_io_ho_input = bc_pe_250_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_251_io_ve_input = bc_pe_219_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_251_io_input_valid = io_input_valid_251; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_251_io_iormac = io_iormac_251; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_252_clock = clock;
  assign bc_pe_252_reset = reset;
  assign bc_pe_252_io_ho_input = bc_pe_251_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_252_io_ve_input = bc_pe_220_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_252_io_input_valid = io_input_valid_252; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_252_io_iormac = io_iormac_252; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_253_clock = clock;
  assign bc_pe_253_reset = reset;
  assign bc_pe_253_io_ho_input = bc_pe_252_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_253_io_ve_input = bc_pe_221_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_253_io_input_valid = io_input_valid_253; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_253_io_iormac = io_iormac_253; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_254_clock = clock;
  assign bc_pe_254_reset = reset;
  assign bc_pe_254_io_ho_input = bc_pe_253_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_254_io_ve_input = bc_pe_222_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_254_io_input_valid = io_input_valid_254; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_254_io_iormac = io_iormac_254; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_255_clock = clock;
  assign bc_pe_255_reset = reset;
  assign bc_pe_255_io_ho_input = bc_pe_254_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_255_io_ve_input = bc_pe_223_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_255_io_input_valid = io_input_valid_255; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_255_io_iormac = io_iormac_255; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_256_clock = clock;
  assign bc_pe_256_reset = reset;
  assign bc_pe_256_io_ho_input = io_x_input_8; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_256_io_ve_input = bc_pe_224_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_256_io_input_valid = io_input_valid_256; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_256_io_iormac = io_iormac_256; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_257_clock = clock;
  assign bc_pe_257_reset = reset;
  assign bc_pe_257_io_ho_input = bc_pe_256_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_257_io_ve_input = bc_pe_225_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_257_io_input_valid = io_input_valid_257; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_257_io_iormac = io_iormac_257; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_258_clock = clock;
  assign bc_pe_258_reset = reset;
  assign bc_pe_258_io_ho_input = bc_pe_257_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_258_io_ve_input = bc_pe_226_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_258_io_input_valid = io_input_valid_258; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_258_io_iormac = io_iormac_258; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_259_clock = clock;
  assign bc_pe_259_reset = reset;
  assign bc_pe_259_io_ho_input = bc_pe_258_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_259_io_ve_input = bc_pe_227_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_259_io_input_valid = io_input_valid_259; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_259_io_iormac = io_iormac_259; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_260_clock = clock;
  assign bc_pe_260_reset = reset;
  assign bc_pe_260_io_ho_input = bc_pe_259_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_260_io_ve_input = bc_pe_228_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_260_io_input_valid = io_input_valid_260; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_260_io_iormac = io_iormac_260; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_261_clock = clock;
  assign bc_pe_261_reset = reset;
  assign bc_pe_261_io_ho_input = bc_pe_260_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_261_io_ve_input = bc_pe_229_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_261_io_input_valid = io_input_valid_261; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_261_io_iormac = io_iormac_261; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_262_clock = clock;
  assign bc_pe_262_reset = reset;
  assign bc_pe_262_io_ho_input = bc_pe_261_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_262_io_ve_input = bc_pe_230_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_262_io_input_valid = io_input_valid_262; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_262_io_iormac = io_iormac_262; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_263_clock = clock;
  assign bc_pe_263_reset = reset;
  assign bc_pe_263_io_ho_input = bc_pe_262_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_263_io_ve_input = bc_pe_231_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_263_io_input_valid = io_input_valid_263; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_263_io_iormac = io_iormac_263; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_264_clock = clock;
  assign bc_pe_264_reset = reset;
  assign bc_pe_264_io_ho_input = bc_pe_263_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_264_io_ve_input = bc_pe_232_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_264_io_input_valid = io_input_valid_264; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_264_io_iormac = io_iormac_264; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_265_clock = clock;
  assign bc_pe_265_reset = reset;
  assign bc_pe_265_io_ho_input = bc_pe_264_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_265_io_ve_input = bc_pe_233_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_265_io_input_valid = io_input_valid_265; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_265_io_iormac = io_iormac_265; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_266_clock = clock;
  assign bc_pe_266_reset = reset;
  assign bc_pe_266_io_ho_input = bc_pe_265_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_266_io_ve_input = bc_pe_234_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_266_io_input_valid = io_input_valid_266; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_266_io_iormac = io_iormac_266; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_267_clock = clock;
  assign bc_pe_267_reset = reset;
  assign bc_pe_267_io_ho_input = bc_pe_266_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_267_io_ve_input = bc_pe_235_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_267_io_input_valid = io_input_valid_267; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_267_io_iormac = io_iormac_267; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_268_clock = clock;
  assign bc_pe_268_reset = reset;
  assign bc_pe_268_io_ho_input = bc_pe_267_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_268_io_ve_input = bc_pe_236_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_268_io_input_valid = io_input_valid_268; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_268_io_iormac = io_iormac_268; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_269_clock = clock;
  assign bc_pe_269_reset = reset;
  assign bc_pe_269_io_ho_input = bc_pe_268_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_269_io_ve_input = bc_pe_237_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_269_io_input_valid = io_input_valid_269; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_269_io_iormac = io_iormac_269; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_270_clock = clock;
  assign bc_pe_270_reset = reset;
  assign bc_pe_270_io_ho_input = bc_pe_269_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_270_io_ve_input = bc_pe_238_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_270_io_input_valid = io_input_valid_270; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_270_io_iormac = io_iormac_270; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_271_clock = clock;
  assign bc_pe_271_reset = reset;
  assign bc_pe_271_io_ho_input = bc_pe_270_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_271_io_ve_input = bc_pe_239_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_271_io_input_valid = io_input_valid_271; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_271_io_iormac = io_iormac_271; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_272_clock = clock;
  assign bc_pe_272_reset = reset;
  assign bc_pe_272_io_ho_input = bc_pe_271_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_272_io_ve_input = bc_pe_240_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_272_io_input_valid = io_input_valid_272; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_272_io_iormac = io_iormac_272; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_273_clock = clock;
  assign bc_pe_273_reset = reset;
  assign bc_pe_273_io_ho_input = bc_pe_272_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_273_io_ve_input = bc_pe_241_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_273_io_input_valid = io_input_valid_273; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_273_io_iormac = io_iormac_273; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_274_clock = clock;
  assign bc_pe_274_reset = reset;
  assign bc_pe_274_io_ho_input = bc_pe_273_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_274_io_ve_input = bc_pe_242_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_274_io_input_valid = io_input_valid_274; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_274_io_iormac = io_iormac_274; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_275_clock = clock;
  assign bc_pe_275_reset = reset;
  assign bc_pe_275_io_ho_input = bc_pe_274_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_275_io_ve_input = bc_pe_243_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_275_io_input_valid = io_input_valid_275; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_275_io_iormac = io_iormac_275; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_276_clock = clock;
  assign bc_pe_276_reset = reset;
  assign bc_pe_276_io_ho_input = bc_pe_275_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_276_io_ve_input = bc_pe_244_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_276_io_input_valid = io_input_valid_276; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_276_io_iormac = io_iormac_276; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_277_clock = clock;
  assign bc_pe_277_reset = reset;
  assign bc_pe_277_io_ho_input = bc_pe_276_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_277_io_ve_input = bc_pe_245_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_277_io_input_valid = io_input_valid_277; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_277_io_iormac = io_iormac_277; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_278_clock = clock;
  assign bc_pe_278_reset = reset;
  assign bc_pe_278_io_ho_input = bc_pe_277_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_278_io_ve_input = bc_pe_246_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_278_io_input_valid = io_input_valid_278; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_278_io_iormac = io_iormac_278; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_279_clock = clock;
  assign bc_pe_279_reset = reset;
  assign bc_pe_279_io_ho_input = bc_pe_278_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_279_io_ve_input = bc_pe_247_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_279_io_input_valid = io_input_valid_279; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_279_io_iormac = io_iormac_279; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_280_clock = clock;
  assign bc_pe_280_reset = reset;
  assign bc_pe_280_io_ho_input = bc_pe_279_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_280_io_ve_input = bc_pe_248_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_280_io_input_valid = io_input_valid_280; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_280_io_iormac = io_iormac_280; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_281_clock = clock;
  assign bc_pe_281_reset = reset;
  assign bc_pe_281_io_ho_input = bc_pe_280_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_281_io_ve_input = bc_pe_249_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_281_io_input_valid = io_input_valid_281; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_281_io_iormac = io_iormac_281; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_282_clock = clock;
  assign bc_pe_282_reset = reset;
  assign bc_pe_282_io_ho_input = bc_pe_281_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_282_io_ve_input = bc_pe_250_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_282_io_input_valid = io_input_valid_282; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_282_io_iormac = io_iormac_282; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_283_clock = clock;
  assign bc_pe_283_reset = reset;
  assign bc_pe_283_io_ho_input = bc_pe_282_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_283_io_ve_input = bc_pe_251_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_283_io_input_valid = io_input_valid_283; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_283_io_iormac = io_iormac_283; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_284_clock = clock;
  assign bc_pe_284_reset = reset;
  assign bc_pe_284_io_ho_input = bc_pe_283_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_284_io_ve_input = bc_pe_252_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_284_io_input_valid = io_input_valid_284; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_284_io_iormac = io_iormac_284; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_285_clock = clock;
  assign bc_pe_285_reset = reset;
  assign bc_pe_285_io_ho_input = bc_pe_284_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_285_io_ve_input = bc_pe_253_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_285_io_input_valid = io_input_valid_285; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_285_io_iormac = io_iormac_285; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_286_clock = clock;
  assign bc_pe_286_reset = reset;
  assign bc_pe_286_io_ho_input = bc_pe_285_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_286_io_ve_input = bc_pe_254_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_286_io_input_valid = io_input_valid_286; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_286_io_iormac = io_iormac_286; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_287_clock = clock;
  assign bc_pe_287_reset = reset;
  assign bc_pe_287_io_ho_input = bc_pe_286_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_287_io_ve_input = bc_pe_255_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_287_io_input_valid = io_input_valid_287; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_287_io_iormac = io_iormac_287; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_288_clock = clock;
  assign bc_pe_288_reset = reset;
  assign bc_pe_288_io_ho_input = io_x_input_9; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_288_io_ve_input = bc_pe_256_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_288_io_input_valid = io_input_valid_288; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_288_io_iormac = io_iormac_288; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_289_clock = clock;
  assign bc_pe_289_reset = reset;
  assign bc_pe_289_io_ho_input = bc_pe_288_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_289_io_ve_input = bc_pe_257_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_289_io_input_valid = io_input_valid_289; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_289_io_iormac = io_iormac_289; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_290_clock = clock;
  assign bc_pe_290_reset = reset;
  assign bc_pe_290_io_ho_input = bc_pe_289_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_290_io_ve_input = bc_pe_258_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_290_io_input_valid = io_input_valid_290; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_290_io_iormac = io_iormac_290; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_291_clock = clock;
  assign bc_pe_291_reset = reset;
  assign bc_pe_291_io_ho_input = bc_pe_290_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_291_io_ve_input = bc_pe_259_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_291_io_input_valid = io_input_valid_291; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_291_io_iormac = io_iormac_291; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_292_clock = clock;
  assign bc_pe_292_reset = reset;
  assign bc_pe_292_io_ho_input = bc_pe_291_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_292_io_ve_input = bc_pe_260_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_292_io_input_valid = io_input_valid_292; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_292_io_iormac = io_iormac_292; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_293_clock = clock;
  assign bc_pe_293_reset = reset;
  assign bc_pe_293_io_ho_input = bc_pe_292_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_293_io_ve_input = bc_pe_261_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_293_io_input_valid = io_input_valid_293; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_293_io_iormac = io_iormac_293; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_294_clock = clock;
  assign bc_pe_294_reset = reset;
  assign bc_pe_294_io_ho_input = bc_pe_293_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_294_io_ve_input = bc_pe_262_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_294_io_input_valid = io_input_valid_294; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_294_io_iormac = io_iormac_294; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_295_clock = clock;
  assign bc_pe_295_reset = reset;
  assign bc_pe_295_io_ho_input = bc_pe_294_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_295_io_ve_input = bc_pe_263_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_295_io_input_valid = io_input_valid_295; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_295_io_iormac = io_iormac_295; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_296_clock = clock;
  assign bc_pe_296_reset = reset;
  assign bc_pe_296_io_ho_input = bc_pe_295_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_296_io_ve_input = bc_pe_264_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_296_io_input_valid = io_input_valid_296; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_296_io_iormac = io_iormac_296; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_297_clock = clock;
  assign bc_pe_297_reset = reset;
  assign bc_pe_297_io_ho_input = bc_pe_296_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_297_io_ve_input = bc_pe_265_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_297_io_input_valid = io_input_valid_297; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_297_io_iormac = io_iormac_297; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_298_clock = clock;
  assign bc_pe_298_reset = reset;
  assign bc_pe_298_io_ho_input = bc_pe_297_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_298_io_ve_input = bc_pe_266_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_298_io_input_valid = io_input_valid_298; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_298_io_iormac = io_iormac_298; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_299_clock = clock;
  assign bc_pe_299_reset = reset;
  assign bc_pe_299_io_ho_input = bc_pe_298_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_299_io_ve_input = bc_pe_267_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_299_io_input_valid = io_input_valid_299; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_299_io_iormac = io_iormac_299; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_300_clock = clock;
  assign bc_pe_300_reset = reset;
  assign bc_pe_300_io_ho_input = bc_pe_299_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_300_io_ve_input = bc_pe_268_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_300_io_input_valid = io_input_valid_300; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_300_io_iormac = io_iormac_300; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_301_clock = clock;
  assign bc_pe_301_reset = reset;
  assign bc_pe_301_io_ho_input = bc_pe_300_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_301_io_ve_input = bc_pe_269_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_301_io_input_valid = io_input_valid_301; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_301_io_iormac = io_iormac_301; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_302_clock = clock;
  assign bc_pe_302_reset = reset;
  assign bc_pe_302_io_ho_input = bc_pe_301_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_302_io_ve_input = bc_pe_270_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_302_io_input_valid = io_input_valid_302; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_302_io_iormac = io_iormac_302; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_303_clock = clock;
  assign bc_pe_303_reset = reset;
  assign bc_pe_303_io_ho_input = bc_pe_302_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_303_io_ve_input = bc_pe_271_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_303_io_input_valid = io_input_valid_303; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_303_io_iormac = io_iormac_303; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_304_clock = clock;
  assign bc_pe_304_reset = reset;
  assign bc_pe_304_io_ho_input = bc_pe_303_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_304_io_ve_input = bc_pe_272_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_304_io_input_valid = io_input_valid_304; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_304_io_iormac = io_iormac_304; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_305_clock = clock;
  assign bc_pe_305_reset = reset;
  assign bc_pe_305_io_ho_input = bc_pe_304_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_305_io_ve_input = bc_pe_273_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_305_io_input_valid = io_input_valid_305; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_305_io_iormac = io_iormac_305; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_306_clock = clock;
  assign bc_pe_306_reset = reset;
  assign bc_pe_306_io_ho_input = bc_pe_305_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_306_io_ve_input = bc_pe_274_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_306_io_input_valid = io_input_valid_306; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_306_io_iormac = io_iormac_306; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_307_clock = clock;
  assign bc_pe_307_reset = reset;
  assign bc_pe_307_io_ho_input = bc_pe_306_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_307_io_ve_input = bc_pe_275_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_307_io_input_valid = io_input_valid_307; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_307_io_iormac = io_iormac_307; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_308_clock = clock;
  assign bc_pe_308_reset = reset;
  assign bc_pe_308_io_ho_input = bc_pe_307_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_308_io_ve_input = bc_pe_276_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_308_io_input_valid = io_input_valid_308; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_308_io_iormac = io_iormac_308; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_309_clock = clock;
  assign bc_pe_309_reset = reset;
  assign bc_pe_309_io_ho_input = bc_pe_308_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_309_io_ve_input = bc_pe_277_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_309_io_input_valid = io_input_valid_309; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_309_io_iormac = io_iormac_309; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_310_clock = clock;
  assign bc_pe_310_reset = reset;
  assign bc_pe_310_io_ho_input = bc_pe_309_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_310_io_ve_input = bc_pe_278_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_310_io_input_valid = io_input_valid_310; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_310_io_iormac = io_iormac_310; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_311_clock = clock;
  assign bc_pe_311_reset = reset;
  assign bc_pe_311_io_ho_input = bc_pe_310_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_311_io_ve_input = bc_pe_279_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_311_io_input_valid = io_input_valid_311; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_311_io_iormac = io_iormac_311; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_312_clock = clock;
  assign bc_pe_312_reset = reset;
  assign bc_pe_312_io_ho_input = bc_pe_311_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_312_io_ve_input = bc_pe_280_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_312_io_input_valid = io_input_valid_312; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_312_io_iormac = io_iormac_312; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_313_clock = clock;
  assign bc_pe_313_reset = reset;
  assign bc_pe_313_io_ho_input = bc_pe_312_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_313_io_ve_input = bc_pe_281_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_313_io_input_valid = io_input_valid_313; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_313_io_iormac = io_iormac_313; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_314_clock = clock;
  assign bc_pe_314_reset = reset;
  assign bc_pe_314_io_ho_input = bc_pe_313_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_314_io_ve_input = bc_pe_282_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_314_io_input_valid = io_input_valid_314; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_314_io_iormac = io_iormac_314; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_315_clock = clock;
  assign bc_pe_315_reset = reset;
  assign bc_pe_315_io_ho_input = bc_pe_314_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_315_io_ve_input = bc_pe_283_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_315_io_input_valid = io_input_valid_315; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_315_io_iormac = io_iormac_315; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_316_clock = clock;
  assign bc_pe_316_reset = reset;
  assign bc_pe_316_io_ho_input = bc_pe_315_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_316_io_ve_input = bc_pe_284_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_316_io_input_valid = io_input_valid_316; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_316_io_iormac = io_iormac_316; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_317_clock = clock;
  assign bc_pe_317_reset = reset;
  assign bc_pe_317_io_ho_input = bc_pe_316_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_317_io_ve_input = bc_pe_285_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_317_io_input_valid = io_input_valid_317; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_317_io_iormac = io_iormac_317; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_318_clock = clock;
  assign bc_pe_318_reset = reset;
  assign bc_pe_318_io_ho_input = bc_pe_317_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_318_io_ve_input = bc_pe_286_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_318_io_input_valid = io_input_valid_318; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_318_io_iormac = io_iormac_318; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_319_clock = clock;
  assign bc_pe_319_reset = reset;
  assign bc_pe_319_io_ho_input = bc_pe_318_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_319_io_ve_input = bc_pe_287_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_319_io_input_valid = io_input_valid_319; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_319_io_iormac = io_iormac_319; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_320_clock = clock;
  assign bc_pe_320_reset = reset;
  assign bc_pe_320_io_ho_input = io_x_input_10; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_320_io_ve_input = bc_pe_288_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_320_io_input_valid = io_input_valid_320; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_320_io_iormac = io_iormac_320; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_321_clock = clock;
  assign bc_pe_321_reset = reset;
  assign bc_pe_321_io_ho_input = bc_pe_320_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_321_io_ve_input = bc_pe_289_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_321_io_input_valid = io_input_valid_321; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_321_io_iormac = io_iormac_321; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_322_clock = clock;
  assign bc_pe_322_reset = reset;
  assign bc_pe_322_io_ho_input = bc_pe_321_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_322_io_ve_input = bc_pe_290_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_322_io_input_valid = io_input_valid_322; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_322_io_iormac = io_iormac_322; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_323_clock = clock;
  assign bc_pe_323_reset = reset;
  assign bc_pe_323_io_ho_input = bc_pe_322_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_323_io_ve_input = bc_pe_291_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_323_io_input_valid = io_input_valid_323; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_323_io_iormac = io_iormac_323; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_324_clock = clock;
  assign bc_pe_324_reset = reset;
  assign bc_pe_324_io_ho_input = bc_pe_323_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_324_io_ve_input = bc_pe_292_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_324_io_input_valid = io_input_valid_324; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_324_io_iormac = io_iormac_324; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_325_clock = clock;
  assign bc_pe_325_reset = reset;
  assign bc_pe_325_io_ho_input = bc_pe_324_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_325_io_ve_input = bc_pe_293_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_325_io_input_valid = io_input_valid_325; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_325_io_iormac = io_iormac_325; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_326_clock = clock;
  assign bc_pe_326_reset = reset;
  assign bc_pe_326_io_ho_input = bc_pe_325_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_326_io_ve_input = bc_pe_294_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_326_io_input_valid = io_input_valid_326; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_326_io_iormac = io_iormac_326; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_327_clock = clock;
  assign bc_pe_327_reset = reset;
  assign bc_pe_327_io_ho_input = bc_pe_326_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_327_io_ve_input = bc_pe_295_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_327_io_input_valid = io_input_valid_327; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_327_io_iormac = io_iormac_327; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_328_clock = clock;
  assign bc_pe_328_reset = reset;
  assign bc_pe_328_io_ho_input = bc_pe_327_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_328_io_ve_input = bc_pe_296_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_328_io_input_valid = io_input_valid_328; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_328_io_iormac = io_iormac_328; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_329_clock = clock;
  assign bc_pe_329_reset = reset;
  assign bc_pe_329_io_ho_input = bc_pe_328_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_329_io_ve_input = bc_pe_297_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_329_io_input_valid = io_input_valid_329; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_329_io_iormac = io_iormac_329; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_330_clock = clock;
  assign bc_pe_330_reset = reset;
  assign bc_pe_330_io_ho_input = bc_pe_329_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_330_io_ve_input = bc_pe_298_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_330_io_input_valid = io_input_valid_330; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_330_io_iormac = io_iormac_330; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_331_clock = clock;
  assign bc_pe_331_reset = reset;
  assign bc_pe_331_io_ho_input = bc_pe_330_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_331_io_ve_input = bc_pe_299_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_331_io_input_valid = io_input_valid_331; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_331_io_iormac = io_iormac_331; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_332_clock = clock;
  assign bc_pe_332_reset = reset;
  assign bc_pe_332_io_ho_input = bc_pe_331_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_332_io_ve_input = bc_pe_300_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_332_io_input_valid = io_input_valid_332; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_332_io_iormac = io_iormac_332; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_333_clock = clock;
  assign bc_pe_333_reset = reset;
  assign bc_pe_333_io_ho_input = bc_pe_332_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_333_io_ve_input = bc_pe_301_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_333_io_input_valid = io_input_valid_333; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_333_io_iormac = io_iormac_333; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_334_clock = clock;
  assign bc_pe_334_reset = reset;
  assign bc_pe_334_io_ho_input = bc_pe_333_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_334_io_ve_input = bc_pe_302_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_334_io_input_valid = io_input_valid_334; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_334_io_iormac = io_iormac_334; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_335_clock = clock;
  assign bc_pe_335_reset = reset;
  assign bc_pe_335_io_ho_input = bc_pe_334_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_335_io_ve_input = bc_pe_303_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_335_io_input_valid = io_input_valid_335; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_335_io_iormac = io_iormac_335; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_336_clock = clock;
  assign bc_pe_336_reset = reset;
  assign bc_pe_336_io_ho_input = bc_pe_335_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_336_io_ve_input = bc_pe_304_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_336_io_input_valid = io_input_valid_336; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_336_io_iormac = io_iormac_336; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_337_clock = clock;
  assign bc_pe_337_reset = reset;
  assign bc_pe_337_io_ho_input = bc_pe_336_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_337_io_ve_input = bc_pe_305_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_337_io_input_valid = io_input_valid_337; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_337_io_iormac = io_iormac_337; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_338_clock = clock;
  assign bc_pe_338_reset = reset;
  assign bc_pe_338_io_ho_input = bc_pe_337_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_338_io_ve_input = bc_pe_306_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_338_io_input_valid = io_input_valid_338; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_338_io_iormac = io_iormac_338; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_339_clock = clock;
  assign bc_pe_339_reset = reset;
  assign bc_pe_339_io_ho_input = bc_pe_338_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_339_io_ve_input = bc_pe_307_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_339_io_input_valid = io_input_valid_339; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_339_io_iormac = io_iormac_339; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_340_clock = clock;
  assign bc_pe_340_reset = reset;
  assign bc_pe_340_io_ho_input = bc_pe_339_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_340_io_ve_input = bc_pe_308_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_340_io_input_valid = io_input_valid_340; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_340_io_iormac = io_iormac_340; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_341_clock = clock;
  assign bc_pe_341_reset = reset;
  assign bc_pe_341_io_ho_input = bc_pe_340_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_341_io_ve_input = bc_pe_309_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_341_io_input_valid = io_input_valid_341; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_341_io_iormac = io_iormac_341; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_342_clock = clock;
  assign bc_pe_342_reset = reset;
  assign bc_pe_342_io_ho_input = bc_pe_341_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_342_io_ve_input = bc_pe_310_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_342_io_input_valid = io_input_valid_342; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_342_io_iormac = io_iormac_342; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_343_clock = clock;
  assign bc_pe_343_reset = reset;
  assign bc_pe_343_io_ho_input = bc_pe_342_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_343_io_ve_input = bc_pe_311_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_343_io_input_valid = io_input_valid_343; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_343_io_iormac = io_iormac_343; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_344_clock = clock;
  assign bc_pe_344_reset = reset;
  assign bc_pe_344_io_ho_input = bc_pe_343_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_344_io_ve_input = bc_pe_312_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_344_io_input_valid = io_input_valid_344; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_344_io_iormac = io_iormac_344; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_345_clock = clock;
  assign bc_pe_345_reset = reset;
  assign bc_pe_345_io_ho_input = bc_pe_344_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_345_io_ve_input = bc_pe_313_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_345_io_input_valid = io_input_valid_345; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_345_io_iormac = io_iormac_345; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_346_clock = clock;
  assign bc_pe_346_reset = reset;
  assign bc_pe_346_io_ho_input = bc_pe_345_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_346_io_ve_input = bc_pe_314_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_346_io_input_valid = io_input_valid_346; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_346_io_iormac = io_iormac_346; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_347_clock = clock;
  assign bc_pe_347_reset = reset;
  assign bc_pe_347_io_ho_input = bc_pe_346_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_347_io_ve_input = bc_pe_315_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_347_io_input_valid = io_input_valid_347; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_347_io_iormac = io_iormac_347; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_348_clock = clock;
  assign bc_pe_348_reset = reset;
  assign bc_pe_348_io_ho_input = bc_pe_347_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_348_io_ve_input = bc_pe_316_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_348_io_input_valid = io_input_valid_348; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_348_io_iormac = io_iormac_348; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_349_clock = clock;
  assign bc_pe_349_reset = reset;
  assign bc_pe_349_io_ho_input = bc_pe_348_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_349_io_ve_input = bc_pe_317_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_349_io_input_valid = io_input_valid_349; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_349_io_iormac = io_iormac_349; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_350_clock = clock;
  assign bc_pe_350_reset = reset;
  assign bc_pe_350_io_ho_input = bc_pe_349_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_350_io_ve_input = bc_pe_318_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_350_io_input_valid = io_input_valid_350; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_350_io_iormac = io_iormac_350; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_351_clock = clock;
  assign bc_pe_351_reset = reset;
  assign bc_pe_351_io_ho_input = bc_pe_350_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_351_io_ve_input = bc_pe_319_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_351_io_input_valid = io_input_valid_351; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_351_io_iormac = io_iormac_351; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_352_clock = clock;
  assign bc_pe_352_reset = reset;
  assign bc_pe_352_io_ho_input = io_x_input_11; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_352_io_ve_input = bc_pe_320_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_352_io_input_valid = io_input_valid_352; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_352_io_iormac = io_iormac_352; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_353_clock = clock;
  assign bc_pe_353_reset = reset;
  assign bc_pe_353_io_ho_input = bc_pe_352_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_353_io_ve_input = bc_pe_321_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_353_io_input_valid = io_input_valid_353; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_353_io_iormac = io_iormac_353; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_354_clock = clock;
  assign bc_pe_354_reset = reset;
  assign bc_pe_354_io_ho_input = bc_pe_353_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_354_io_ve_input = bc_pe_322_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_354_io_input_valid = io_input_valid_354; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_354_io_iormac = io_iormac_354; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_355_clock = clock;
  assign bc_pe_355_reset = reset;
  assign bc_pe_355_io_ho_input = bc_pe_354_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_355_io_ve_input = bc_pe_323_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_355_io_input_valid = io_input_valid_355; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_355_io_iormac = io_iormac_355; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_356_clock = clock;
  assign bc_pe_356_reset = reset;
  assign bc_pe_356_io_ho_input = bc_pe_355_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_356_io_ve_input = bc_pe_324_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_356_io_input_valid = io_input_valid_356; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_356_io_iormac = io_iormac_356; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_357_clock = clock;
  assign bc_pe_357_reset = reset;
  assign bc_pe_357_io_ho_input = bc_pe_356_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_357_io_ve_input = bc_pe_325_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_357_io_input_valid = io_input_valid_357; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_357_io_iormac = io_iormac_357; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_358_clock = clock;
  assign bc_pe_358_reset = reset;
  assign bc_pe_358_io_ho_input = bc_pe_357_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_358_io_ve_input = bc_pe_326_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_358_io_input_valid = io_input_valid_358; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_358_io_iormac = io_iormac_358; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_359_clock = clock;
  assign bc_pe_359_reset = reset;
  assign bc_pe_359_io_ho_input = bc_pe_358_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_359_io_ve_input = bc_pe_327_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_359_io_input_valid = io_input_valid_359; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_359_io_iormac = io_iormac_359; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_360_clock = clock;
  assign bc_pe_360_reset = reset;
  assign bc_pe_360_io_ho_input = bc_pe_359_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_360_io_ve_input = bc_pe_328_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_360_io_input_valid = io_input_valid_360; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_360_io_iormac = io_iormac_360; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_361_clock = clock;
  assign bc_pe_361_reset = reset;
  assign bc_pe_361_io_ho_input = bc_pe_360_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_361_io_ve_input = bc_pe_329_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_361_io_input_valid = io_input_valid_361; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_361_io_iormac = io_iormac_361; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_362_clock = clock;
  assign bc_pe_362_reset = reset;
  assign bc_pe_362_io_ho_input = bc_pe_361_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_362_io_ve_input = bc_pe_330_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_362_io_input_valid = io_input_valid_362; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_362_io_iormac = io_iormac_362; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_363_clock = clock;
  assign bc_pe_363_reset = reset;
  assign bc_pe_363_io_ho_input = bc_pe_362_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_363_io_ve_input = bc_pe_331_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_363_io_input_valid = io_input_valid_363; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_363_io_iormac = io_iormac_363; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_364_clock = clock;
  assign bc_pe_364_reset = reset;
  assign bc_pe_364_io_ho_input = bc_pe_363_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_364_io_ve_input = bc_pe_332_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_364_io_input_valid = io_input_valid_364; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_364_io_iormac = io_iormac_364; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_365_clock = clock;
  assign bc_pe_365_reset = reset;
  assign bc_pe_365_io_ho_input = bc_pe_364_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_365_io_ve_input = bc_pe_333_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_365_io_input_valid = io_input_valid_365; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_365_io_iormac = io_iormac_365; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_366_clock = clock;
  assign bc_pe_366_reset = reset;
  assign bc_pe_366_io_ho_input = bc_pe_365_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_366_io_ve_input = bc_pe_334_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_366_io_input_valid = io_input_valid_366; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_366_io_iormac = io_iormac_366; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_367_clock = clock;
  assign bc_pe_367_reset = reset;
  assign bc_pe_367_io_ho_input = bc_pe_366_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_367_io_ve_input = bc_pe_335_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_367_io_input_valid = io_input_valid_367; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_367_io_iormac = io_iormac_367; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_368_clock = clock;
  assign bc_pe_368_reset = reset;
  assign bc_pe_368_io_ho_input = bc_pe_367_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_368_io_ve_input = bc_pe_336_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_368_io_input_valid = io_input_valid_368; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_368_io_iormac = io_iormac_368; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_369_clock = clock;
  assign bc_pe_369_reset = reset;
  assign bc_pe_369_io_ho_input = bc_pe_368_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_369_io_ve_input = bc_pe_337_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_369_io_input_valid = io_input_valid_369; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_369_io_iormac = io_iormac_369; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_370_clock = clock;
  assign bc_pe_370_reset = reset;
  assign bc_pe_370_io_ho_input = bc_pe_369_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_370_io_ve_input = bc_pe_338_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_370_io_input_valid = io_input_valid_370; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_370_io_iormac = io_iormac_370; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_371_clock = clock;
  assign bc_pe_371_reset = reset;
  assign bc_pe_371_io_ho_input = bc_pe_370_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_371_io_ve_input = bc_pe_339_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_371_io_input_valid = io_input_valid_371; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_371_io_iormac = io_iormac_371; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_372_clock = clock;
  assign bc_pe_372_reset = reset;
  assign bc_pe_372_io_ho_input = bc_pe_371_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_372_io_ve_input = bc_pe_340_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_372_io_input_valid = io_input_valid_372; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_372_io_iormac = io_iormac_372; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_373_clock = clock;
  assign bc_pe_373_reset = reset;
  assign bc_pe_373_io_ho_input = bc_pe_372_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_373_io_ve_input = bc_pe_341_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_373_io_input_valid = io_input_valid_373; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_373_io_iormac = io_iormac_373; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_374_clock = clock;
  assign bc_pe_374_reset = reset;
  assign bc_pe_374_io_ho_input = bc_pe_373_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_374_io_ve_input = bc_pe_342_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_374_io_input_valid = io_input_valid_374; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_374_io_iormac = io_iormac_374; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_375_clock = clock;
  assign bc_pe_375_reset = reset;
  assign bc_pe_375_io_ho_input = bc_pe_374_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_375_io_ve_input = bc_pe_343_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_375_io_input_valid = io_input_valid_375; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_375_io_iormac = io_iormac_375; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_376_clock = clock;
  assign bc_pe_376_reset = reset;
  assign bc_pe_376_io_ho_input = bc_pe_375_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_376_io_ve_input = bc_pe_344_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_376_io_input_valid = io_input_valid_376; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_376_io_iormac = io_iormac_376; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_377_clock = clock;
  assign bc_pe_377_reset = reset;
  assign bc_pe_377_io_ho_input = bc_pe_376_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_377_io_ve_input = bc_pe_345_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_377_io_input_valid = io_input_valid_377; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_377_io_iormac = io_iormac_377; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_378_clock = clock;
  assign bc_pe_378_reset = reset;
  assign bc_pe_378_io_ho_input = bc_pe_377_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_378_io_ve_input = bc_pe_346_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_378_io_input_valid = io_input_valid_378; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_378_io_iormac = io_iormac_378; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_379_clock = clock;
  assign bc_pe_379_reset = reset;
  assign bc_pe_379_io_ho_input = bc_pe_378_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_379_io_ve_input = bc_pe_347_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_379_io_input_valid = io_input_valid_379; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_379_io_iormac = io_iormac_379; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_380_clock = clock;
  assign bc_pe_380_reset = reset;
  assign bc_pe_380_io_ho_input = bc_pe_379_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_380_io_ve_input = bc_pe_348_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_380_io_input_valid = io_input_valid_380; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_380_io_iormac = io_iormac_380; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_381_clock = clock;
  assign bc_pe_381_reset = reset;
  assign bc_pe_381_io_ho_input = bc_pe_380_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_381_io_ve_input = bc_pe_349_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_381_io_input_valid = io_input_valid_381; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_381_io_iormac = io_iormac_381; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_382_clock = clock;
  assign bc_pe_382_reset = reset;
  assign bc_pe_382_io_ho_input = bc_pe_381_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_382_io_ve_input = bc_pe_350_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_382_io_input_valid = io_input_valid_382; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_382_io_iormac = io_iormac_382; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_383_clock = clock;
  assign bc_pe_383_reset = reset;
  assign bc_pe_383_io_ho_input = bc_pe_382_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_383_io_ve_input = bc_pe_351_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_383_io_input_valid = io_input_valid_383; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_383_io_iormac = io_iormac_383; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_384_clock = clock;
  assign bc_pe_384_reset = reset;
  assign bc_pe_384_io_ho_input = io_x_input_12; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_384_io_ve_input = bc_pe_352_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_384_io_input_valid = io_input_valid_384; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_384_io_iormac = io_iormac_384; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_385_clock = clock;
  assign bc_pe_385_reset = reset;
  assign bc_pe_385_io_ho_input = bc_pe_384_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_385_io_ve_input = bc_pe_353_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_385_io_input_valid = io_input_valid_385; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_385_io_iormac = io_iormac_385; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_386_clock = clock;
  assign bc_pe_386_reset = reset;
  assign bc_pe_386_io_ho_input = bc_pe_385_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_386_io_ve_input = bc_pe_354_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_386_io_input_valid = io_input_valid_386; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_386_io_iormac = io_iormac_386; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_387_clock = clock;
  assign bc_pe_387_reset = reset;
  assign bc_pe_387_io_ho_input = bc_pe_386_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_387_io_ve_input = bc_pe_355_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_387_io_input_valid = io_input_valid_387; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_387_io_iormac = io_iormac_387; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_388_clock = clock;
  assign bc_pe_388_reset = reset;
  assign bc_pe_388_io_ho_input = bc_pe_387_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_388_io_ve_input = bc_pe_356_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_388_io_input_valid = io_input_valid_388; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_388_io_iormac = io_iormac_388; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_389_clock = clock;
  assign bc_pe_389_reset = reset;
  assign bc_pe_389_io_ho_input = bc_pe_388_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_389_io_ve_input = bc_pe_357_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_389_io_input_valid = io_input_valid_389; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_389_io_iormac = io_iormac_389; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_390_clock = clock;
  assign bc_pe_390_reset = reset;
  assign bc_pe_390_io_ho_input = bc_pe_389_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_390_io_ve_input = bc_pe_358_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_390_io_input_valid = io_input_valid_390; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_390_io_iormac = io_iormac_390; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_391_clock = clock;
  assign bc_pe_391_reset = reset;
  assign bc_pe_391_io_ho_input = bc_pe_390_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_391_io_ve_input = bc_pe_359_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_391_io_input_valid = io_input_valid_391; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_391_io_iormac = io_iormac_391; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_392_clock = clock;
  assign bc_pe_392_reset = reset;
  assign bc_pe_392_io_ho_input = bc_pe_391_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_392_io_ve_input = bc_pe_360_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_392_io_input_valid = io_input_valid_392; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_392_io_iormac = io_iormac_392; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_393_clock = clock;
  assign bc_pe_393_reset = reset;
  assign bc_pe_393_io_ho_input = bc_pe_392_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_393_io_ve_input = bc_pe_361_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_393_io_input_valid = io_input_valid_393; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_393_io_iormac = io_iormac_393; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_394_clock = clock;
  assign bc_pe_394_reset = reset;
  assign bc_pe_394_io_ho_input = bc_pe_393_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_394_io_ve_input = bc_pe_362_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_394_io_input_valid = io_input_valid_394; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_394_io_iormac = io_iormac_394; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_395_clock = clock;
  assign bc_pe_395_reset = reset;
  assign bc_pe_395_io_ho_input = bc_pe_394_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_395_io_ve_input = bc_pe_363_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_395_io_input_valid = io_input_valid_395; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_395_io_iormac = io_iormac_395; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_396_clock = clock;
  assign bc_pe_396_reset = reset;
  assign bc_pe_396_io_ho_input = bc_pe_395_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_396_io_ve_input = bc_pe_364_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_396_io_input_valid = io_input_valid_396; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_396_io_iormac = io_iormac_396; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_397_clock = clock;
  assign bc_pe_397_reset = reset;
  assign bc_pe_397_io_ho_input = bc_pe_396_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_397_io_ve_input = bc_pe_365_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_397_io_input_valid = io_input_valid_397; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_397_io_iormac = io_iormac_397; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_398_clock = clock;
  assign bc_pe_398_reset = reset;
  assign bc_pe_398_io_ho_input = bc_pe_397_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_398_io_ve_input = bc_pe_366_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_398_io_input_valid = io_input_valid_398; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_398_io_iormac = io_iormac_398; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_399_clock = clock;
  assign bc_pe_399_reset = reset;
  assign bc_pe_399_io_ho_input = bc_pe_398_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_399_io_ve_input = bc_pe_367_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_399_io_input_valid = io_input_valid_399; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_399_io_iormac = io_iormac_399; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_400_clock = clock;
  assign bc_pe_400_reset = reset;
  assign bc_pe_400_io_ho_input = bc_pe_399_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_400_io_ve_input = bc_pe_368_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_400_io_input_valid = io_input_valid_400; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_400_io_iormac = io_iormac_400; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_401_clock = clock;
  assign bc_pe_401_reset = reset;
  assign bc_pe_401_io_ho_input = bc_pe_400_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_401_io_ve_input = bc_pe_369_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_401_io_input_valid = io_input_valid_401; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_401_io_iormac = io_iormac_401; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_402_clock = clock;
  assign bc_pe_402_reset = reset;
  assign bc_pe_402_io_ho_input = bc_pe_401_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_402_io_ve_input = bc_pe_370_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_402_io_input_valid = io_input_valid_402; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_402_io_iormac = io_iormac_402; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_403_clock = clock;
  assign bc_pe_403_reset = reset;
  assign bc_pe_403_io_ho_input = bc_pe_402_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_403_io_ve_input = bc_pe_371_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_403_io_input_valid = io_input_valid_403; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_403_io_iormac = io_iormac_403; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_404_clock = clock;
  assign bc_pe_404_reset = reset;
  assign bc_pe_404_io_ho_input = bc_pe_403_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_404_io_ve_input = bc_pe_372_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_404_io_input_valid = io_input_valid_404; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_404_io_iormac = io_iormac_404; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_405_clock = clock;
  assign bc_pe_405_reset = reset;
  assign bc_pe_405_io_ho_input = bc_pe_404_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_405_io_ve_input = bc_pe_373_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_405_io_input_valid = io_input_valid_405; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_405_io_iormac = io_iormac_405; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_406_clock = clock;
  assign bc_pe_406_reset = reset;
  assign bc_pe_406_io_ho_input = bc_pe_405_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_406_io_ve_input = bc_pe_374_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_406_io_input_valid = io_input_valid_406; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_406_io_iormac = io_iormac_406; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_407_clock = clock;
  assign bc_pe_407_reset = reset;
  assign bc_pe_407_io_ho_input = bc_pe_406_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_407_io_ve_input = bc_pe_375_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_407_io_input_valid = io_input_valid_407; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_407_io_iormac = io_iormac_407; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_408_clock = clock;
  assign bc_pe_408_reset = reset;
  assign bc_pe_408_io_ho_input = bc_pe_407_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_408_io_ve_input = bc_pe_376_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_408_io_input_valid = io_input_valid_408; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_408_io_iormac = io_iormac_408; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_409_clock = clock;
  assign bc_pe_409_reset = reset;
  assign bc_pe_409_io_ho_input = bc_pe_408_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_409_io_ve_input = bc_pe_377_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_409_io_input_valid = io_input_valid_409; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_409_io_iormac = io_iormac_409; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_410_clock = clock;
  assign bc_pe_410_reset = reset;
  assign bc_pe_410_io_ho_input = bc_pe_409_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_410_io_ve_input = bc_pe_378_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_410_io_input_valid = io_input_valid_410; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_410_io_iormac = io_iormac_410; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_411_clock = clock;
  assign bc_pe_411_reset = reset;
  assign bc_pe_411_io_ho_input = bc_pe_410_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_411_io_ve_input = bc_pe_379_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_411_io_input_valid = io_input_valid_411; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_411_io_iormac = io_iormac_411; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_412_clock = clock;
  assign bc_pe_412_reset = reset;
  assign bc_pe_412_io_ho_input = bc_pe_411_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_412_io_ve_input = bc_pe_380_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_412_io_input_valid = io_input_valid_412; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_412_io_iormac = io_iormac_412; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_413_clock = clock;
  assign bc_pe_413_reset = reset;
  assign bc_pe_413_io_ho_input = bc_pe_412_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_413_io_ve_input = bc_pe_381_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_413_io_input_valid = io_input_valid_413; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_413_io_iormac = io_iormac_413; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_414_clock = clock;
  assign bc_pe_414_reset = reset;
  assign bc_pe_414_io_ho_input = bc_pe_413_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_414_io_ve_input = bc_pe_382_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_414_io_input_valid = io_input_valid_414; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_414_io_iormac = io_iormac_414; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_415_clock = clock;
  assign bc_pe_415_reset = reset;
  assign bc_pe_415_io_ho_input = bc_pe_414_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_415_io_ve_input = bc_pe_383_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_415_io_input_valid = io_input_valid_415; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_415_io_iormac = io_iormac_415; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_416_clock = clock;
  assign bc_pe_416_reset = reset;
  assign bc_pe_416_io_ho_input = io_x_input_13; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_416_io_ve_input = bc_pe_384_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_416_io_input_valid = io_input_valid_416; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_416_io_iormac = io_iormac_416; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_417_clock = clock;
  assign bc_pe_417_reset = reset;
  assign bc_pe_417_io_ho_input = bc_pe_416_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_417_io_ve_input = bc_pe_385_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_417_io_input_valid = io_input_valid_417; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_417_io_iormac = io_iormac_417; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_418_clock = clock;
  assign bc_pe_418_reset = reset;
  assign bc_pe_418_io_ho_input = bc_pe_417_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_418_io_ve_input = bc_pe_386_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_418_io_input_valid = io_input_valid_418; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_418_io_iormac = io_iormac_418; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_419_clock = clock;
  assign bc_pe_419_reset = reset;
  assign bc_pe_419_io_ho_input = bc_pe_418_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_419_io_ve_input = bc_pe_387_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_419_io_input_valid = io_input_valid_419; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_419_io_iormac = io_iormac_419; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_420_clock = clock;
  assign bc_pe_420_reset = reset;
  assign bc_pe_420_io_ho_input = bc_pe_419_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_420_io_ve_input = bc_pe_388_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_420_io_input_valid = io_input_valid_420; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_420_io_iormac = io_iormac_420; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_421_clock = clock;
  assign bc_pe_421_reset = reset;
  assign bc_pe_421_io_ho_input = bc_pe_420_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_421_io_ve_input = bc_pe_389_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_421_io_input_valid = io_input_valid_421; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_421_io_iormac = io_iormac_421; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_422_clock = clock;
  assign bc_pe_422_reset = reset;
  assign bc_pe_422_io_ho_input = bc_pe_421_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_422_io_ve_input = bc_pe_390_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_422_io_input_valid = io_input_valid_422; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_422_io_iormac = io_iormac_422; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_423_clock = clock;
  assign bc_pe_423_reset = reset;
  assign bc_pe_423_io_ho_input = bc_pe_422_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_423_io_ve_input = bc_pe_391_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_423_io_input_valid = io_input_valid_423; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_423_io_iormac = io_iormac_423; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_424_clock = clock;
  assign bc_pe_424_reset = reset;
  assign bc_pe_424_io_ho_input = bc_pe_423_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_424_io_ve_input = bc_pe_392_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_424_io_input_valid = io_input_valid_424; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_424_io_iormac = io_iormac_424; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_425_clock = clock;
  assign bc_pe_425_reset = reset;
  assign bc_pe_425_io_ho_input = bc_pe_424_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_425_io_ve_input = bc_pe_393_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_425_io_input_valid = io_input_valid_425; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_425_io_iormac = io_iormac_425; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_426_clock = clock;
  assign bc_pe_426_reset = reset;
  assign bc_pe_426_io_ho_input = bc_pe_425_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_426_io_ve_input = bc_pe_394_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_426_io_input_valid = io_input_valid_426; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_426_io_iormac = io_iormac_426; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_427_clock = clock;
  assign bc_pe_427_reset = reset;
  assign bc_pe_427_io_ho_input = bc_pe_426_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_427_io_ve_input = bc_pe_395_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_427_io_input_valid = io_input_valid_427; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_427_io_iormac = io_iormac_427; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_428_clock = clock;
  assign bc_pe_428_reset = reset;
  assign bc_pe_428_io_ho_input = bc_pe_427_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_428_io_ve_input = bc_pe_396_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_428_io_input_valid = io_input_valid_428; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_428_io_iormac = io_iormac_428; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_429_clock = clock;
  assign bc_pe_429_reset = reset;
  assign bc_pe_429_io_ho_input = bc_pe_428_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_429_io_ve_input = bc_pe_397_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_429_io_input_valid = io_input_valid_429; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_429_io_iormac = io_iormac_429; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_430_clock = clock;
  assign bc_pe_430_reset = reset;
  assign bc_pe_430_io_ho_input = bc_pe_429_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_430_io_ve_input = bc_pe_398_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_430_io_input_valid = io_input_valid_430; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_430_io_iormac = io_iormac_430; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_431_clock = clock;
  assign bc_pe_431_reset = reset;
  assign bc_pe_431_io_ho_input = bc_pe_430_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_431_io_ve_input = bc_pe_399_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_431_io_input_valid = io_input_valid_431; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_431_io_iormac = io_iormac_431; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_432_clock = clock;
  assign bc_pe_432_reset = reset;
  assign bc_pe_432_io_ho_input = bc_pe_431_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_432_io_ve_input = bc_pe_400_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_432_io_input_valid = io_input_valid_432; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_432_io_iormac = io_iormac_432; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_433_clock = clock;
  assign bc_pe_433_reset = reset;
  assign bc_pe_433_io_ho_input = bc_pe_432_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_433_io_ve_input = bc_pe_401_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_433_io_input_valid = io_input_valid_433; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_433_io_iormac = io_iormac_433; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_434_clock = clock;
  assign bc_pe_434_reset = reset;
  assign bc_pe_434_io_ho_input = bc_pe_433_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_434_io_ve_input = bc_pe_402_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_434_io_input_valid = io_input_valid_434; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_434_io_iormac = io_iormac_434; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_435_clock = clock;
  assign bc_pe_435_reset = reset;
  assign bc_pe_435_io_ho_input = bc_pe_434_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_435_io_ve_input = bc_pe_403_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_435_io_input_valid = io_input_valid_435; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_435_io_iormac = io_iormac_435; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_436_clock = clock;
  assign bc_pe_436_reset = reset;
  assign bc_pe_436_io_ho_input = bc_pe_435_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_436_io_ve_input = bc_pe_404_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_436_io_input_valid = io_input_valid_436; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_436_io_iormac = io_iormac_436; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_437_clock = clock;
  assign bc_pe_437_reset = reset;
  assign bc_pe_437_io_ho_input = bc_pe_436_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_437_io_ve_input = bc_pe_405_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_437_io_input_valid = io_input_valid_437; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_437_io_iormac = io_iormac_437; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_438_clock = clock;
  assign bc_pe_438_reset = reset;
  assign bc_pe_438_io_ho_input = bc_pe_437_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_438_io_ve_input = bc_pe_406_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_438_io_input_valid = io_input_valid_438; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_438_io_iormac = io_iormac_438; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_439_clock = clock;
  assign bc_pe_439_reset = reset;
  assign bc_pe_439_io_ho_input = bc_pe_438_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_439_io_ve_input = bc_pe_407_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_439_io_input_valid = io_input_valid_439; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_439_io_iormac = io_iormac_439; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_440_clock = clock;
  assign bc_pe_440_reset = reset;
  assign bc_pe_440_io_ho_input = bc_pe_439_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_440_io_ve_input = bc_pe_408_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_440_io_input_valid = io_input_valid_440; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_440_io_iormac = io_iormac_440; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_441_clock = clock;
  assign bc_pe_441_reset = reset;
  assign bc_pe_441_io_ho_input = bc_pe_440_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_441_io_ve_input = bc_pe_409_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_441_io_input_valid = io_input_valid_441; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_441_io_iormac = io_iormac_441; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_442_clock = clock;
  assign bc_pe_442_reset = reset;
  assign bc_pe_442_io_ho_input = bc_pe_441_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_442_io_ve_input = bc_pe_410_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_442_io_input_valid = io_input_valid_442; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_442_io_iormac = io_iormac_442; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_443_clock = clock;
  assign bc_pe_443_reset = reset;
  assign bc_pe_443_io_ho_input = bc_pe_442_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_443_io_ve_input = bc_pe_411_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_443_io_input_valid = io_input_valid_443; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_443_io_iormac = io_iormac_443; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_444_clock = clock;
  assign bc_pe_444_reset = reset;
  assign bc_pe_444_io_ho_input = bc_pe_443_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_444_io_ve_input = bc_pe_412_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_444_io_input_valid = io_input_valid_444; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_444_io_iormac = io_iormac_444; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_445_clock = clock;
  assign bc_pe_445_reset = reset;
  assign bc_pe_445_io_ho_input = bc_pe_444_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_445_io_ve_input = bc_pe_413_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_445_io_input_valid = io_input_valid_445; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_445_io_iormac = io_iormac_445; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_446_clock = clock;
  assign bc_pe_446_reset = reset;
  assign bc_pe_446_io_ho_input = bc_pe_445_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_446_io_ve_input = bc_pe_414_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_446_io_input_valid = io_input_valid_446; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_446_io_iormac = io_iormac_446; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_447_clock = clock;
  assign bc_pe_447_reset = reset;
  assign bc_pe_447_io_ho_input = bc_pe_446_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_447_io_ve_input = bc_pe_415_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_447_io_input_valid = io_input_valid_447; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_447_io_iormac = io_iormac_447; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_448_clock = clock;
  assign bc_pe_448_reset = reset;
  assign bc_pe_448_io_ho_input = io_x_input_14; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_448_io_ve_input = bc_pe_416_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_448_io_input_valid = io_input_valid_448; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_448_io_iormac = io_iormac_448; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_449_clock = clock;
  assign bc_pe_449_reset = reset;
  assign bc_pe_449_io_ho_input = bc_pe_448_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_449_io_ve_input = bc_pe_417_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_449_io_input_valid = io_input_valid_449; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_449_io_iormac = io_iormac_449; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_450_clock = clock;
  assign bc_pe_450_reset = reset;
  assign bc_pe_450_io_ho_input = bc_pe_449_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_450_io_ve_input = bc_pe_418_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_450_io_input_valid = io_input_valid_450; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_450_io_iormac = io_iormac_450; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_451_clock = clock;
  assign bc_pe_451_reset = reset;
  assign bc_pe_451_io_ho_input = bc_pe_450_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_451_io_ve_input = bc_pe_419_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_451_io_input_valid = io_input_valid_451; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_451_io_iormac = io_iormac_451; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_452_clock = clock;
  assign bc_pe_452_reset = reset;
  assign bc_pe_452_io_ho_input = bc_pe_451_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_452_io_ve_input = bc_pe_420_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_452_io_input_valid = io_input_valid_452; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_452_io_iormac = io_iormac_452; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_453_clock = clock;
  assign bc_pe_453_reset = reset;
  assign bc_pe_453_io_ho_input = bc_pe_452_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_453_io_ve_input = bc_pe_421_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_453_io_input_valid = io_input_valid_453; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_453_io_iormac = io_iormac_453; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_454_clock = clock;
  assign bc_pe_454_reset = reset;
  assign bc_pe_454_io_ho_input = bc_pe_453_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_454_io_ve_input = bc_pe_422_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_454_io_input_valid = io_input_valid_454; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_454_io_iormac = io_iormac_454; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_455_clock = clock;
  assign bc_pe_455_reset = reset;
  assign bc_pe_455_io_ho_input = bc_pe_454_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_455_io_ve_input = bc_pe_423_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_455_io_input_valid = io_input_valid_455; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_455_io_iormac = io_iormac_455; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_456_clock = clock;
  assign bc_pe_456_reset = reset;
  assign bc_pe_456_io_ho_input = bc_pe_455_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_456_io_ve_input = bc_pe_424_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_456_io_input_valid = io_input_valid_456; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_456_io_iormac = io_iormac_456; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_457_clock = clock;
  assign bc_pe_457_reset = reset;
  assign bc_pe_457_io_ho_input = bc_pe_456_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_457_io_ve_input = bc_pe_425_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_457_io_input_valid = io_input_valid_457; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_457_io_iormac = io_iormac_457; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_458_clock = clock;
  assign bc_pe_458_reset = reset;
  assign bc_pe_458_io_ho_input = bc_pe_457_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_458_io_ve_input = bc_pe_426_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_458_io_input_valid = io_input_valid_458; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_458_io_iormac = io_iormac_458; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_459_clock = clock;
  assign bc_pe_459_reset = reset;
  assign bc_pe_459_io_ho_input = bc_pe_458_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_459_io_ve_input = bc_pe_427_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_459_io_input_valid = io_input_valid_459; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_459_io_iormac = io_iormac_459; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_460_clock = clock;
  assign bc_pe_460_reset = reset;
  assign bc_pe_460_io_ho_input = bc_pe_459_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_460_io_ve_input = bc_pe_428_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_460_io_input_valid = io_input_valid_460; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_460_io_iormac = io_iormac_460; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_461_clock = clock;
  assign bc_pe_461_reset = reset;
  assign bc_pe_461_io_ho_input = bc_pe_460_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_461_io_ve_input = bc_pe_429_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_461_io_input_valid = io_input_valid_461; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_461_io_iormac = io_iormac_461; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_462_clock = clock;
  assign bc_pe_462_reset = reset;
  assign bc_pe_462_io_ho_input = bc_pe_461_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_462_io_ve_input = bc_pe_430_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_462_io_input_valid = io_input_valid_462; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_462_io_iormac = io_iormac_462; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_463_clock = clock;
  assign bc_pe_463_reset = reset;
  assign bc_pe_463_io_ho_input = bc_pe_462_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_463_io_ve_input = bc_pe_431_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_463_io_input_valid = io_input_valid_463; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_463_io_iormac = io_iormac_463; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_464_clock = clock;
  assign bc_pe_464_reset = reset;
  assign bc_pe_464_io_ho_input = bc_pe_463_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_464_io_ve_input = bc_pe_432_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_464_io_input_valid = io_input_valid_464; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_464_io_iormac = io_iormac_464; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_465_clock = clock;
  assign bc_pe_465_reset = reset;
  assign bc_pe_465_io_ho_input = bc_pe_464_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_465_io_ve_input = bc_pe_433_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_465_io_input_valid = io_input_valid_465; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_465_io_iormac = io_iormac_465; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_466_clock = clock;
  assign bc_pe_466_reset = reset;
  assign bc_pe_466_io_ho_input = bc_pe_465_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_466_io_ve_input = bc_pe_434_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_466_io_input_valid = io_input_valid_466; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_466_io_iormac = io_iormac_466; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_467_clock = clock;
  assign bc_pe_467_reset = reset;
  assign bc_pe_467_io_ho_input = bc_pe_466_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_467_io_ve_input = bc_pe_435_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_467_io_input_valid = io_input_valid_467; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_467_io_iormac = io_iormac_467; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_468_clock = clock;
  assign bc_pe_468_reset = reset;
  assign bc_pe_468_io_ho_input = bc_pe_467_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_468_io_ve_input = bc_pe_436_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_468_io_input_valid = io_input_valid_468; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_468_io_iormac = io_iormac_468; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_469_clock = clock;
  assign bc_pe_469_reset = reset;
  assign bc_pe_469_io_ho_input = bc_pe_468_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_469_io_ve_input = bc_pe_437_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_469_io_input_valid = io_input_valid_469; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_469_io_iormac = io_iormac_469; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_470_clock = clock;
  assign bc_pe_470_reset = reset;
  assign bc_pe_470_io_ho_input = bc_pe_469_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_470_io_ve_input = bc_pe_438_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_470_io_input_valid = io_input_valid_470; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_470_io_iormac = io_iormac_470; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_471_clock = clock;
  assign bc_pe_471_reset = reset;
  assign bc_pe_471_io_ho_input = bc_pe_470_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_471_io_ve_input = bc_pe_439_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_471_io_input_valid = io_input_valid_471; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_471_io_iormac = io_iormac_471; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_472_clock = clock;
  assign bc_pe_472_reset = reset;
  assign bc_pe_472_io_ho_input = bc_pe_471_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_472_io_ve_input = bc_pe_440_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_472_io_input_valid = io_input_valid_472; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_472_io_iormac = io_iormac_472; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_473_clock = clock;
  assign bc_pe_473_reset = reset;
  assign bc_pe_473_io_ho_input = bc_pe_472_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_473_io_ve_input = bc_pe_441_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_473_io_input_valid = io_input_valid_473; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_473_io_iormac = io_iormac_473; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_474_clock = clock;
  assign bc_pe_474_reset = reset;
  assign bc_pe_474_io_ho_input = bc_pe_473_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_474_io_ve_input = bc_pe_442_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_474_io_input_valid = io_input_valid_474; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_474_io_iormac = io_iormac_474; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_475_clock = clock;
  assign bc_pe_475_reset = reset;
  assign bc_pe_475_io_ho_input = bc_pe_474_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_475_io_ve_input = bc_pe_443_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_475_io_input_valid = io_input_valid_475; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_475_io_iormac = io_iormac_475; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_476_clock = clock;
  assign bc_pe_476_reset = reset;
  assign bc_pe_476_io_ho_input = bc_pe_475_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_476_io_ve_input = bc_pe_444_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_476_io_input_valid = io_input_valid_476; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_476_io_iormac = io_iormac_476; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_477_clock = clock;
  assign bc_pe_477_reset = reset;
  assign bc_pe_477_io_ho_input = bc_pe_476_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_477_io_ve_input = bc_pe_445_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_477_io_input_valid = io_input_valid_477; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_477_io_iormac = io_iormac_477; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_478_clock = clock;
  assign bc_pe_478_reset = reset;
  assign bc_pe_478_io_ho_input = bc_pe_477_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_478_io_ve_input = bc_pe_446_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_478_io_input_valid = io_input_valid_478; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_478_io_iormac = io_iormac_478; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_479_clock = clock;
  assign bc_pe_479_reset = reset;
  assign bc_pe_479_io_ho_input = bc_pe_478_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_479_io_ve_input = bc_pe_447_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_479_io_input_valid = io_input_valid_479; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_479_io_iormac = io_iormac_479; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_480_clock = clock;
  assign bc_pe_480_reset = reset;
  assign bc_pe_480_io_ho_input = io_x_input_15; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_480_io_ve_input = bc_pe_448_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_480_io_input_valid = io_input_valid_480; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_480_io_iormac = io_iormac_480; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_481_clock = clock;
  assign bc_pe_481_reset = reset;
  assign bc_pe_481_io_ho_input = bc_pe_480_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_481_io_ve_input = bc_pe_449_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_481_io_input_valid = io_input_valid_481; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_481_io_iormac = io_iormac_481; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_482_clock = clock;
  assign bc_pe_482_reset = reset;
  assign bc_pe_482_io_ho_input = bc_pe_481_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_482_io_ve_input = bc_pe_450_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_482_io_input_valid = io_input_valid_482; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_482_io_iormac = io_iormac_482; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_483_clock = clock;
  assign bc_pe_483_reset = reset;
  assign bc_pe_483_io_ho_input = bc_pe_482_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_483_io_ve_input = bc_pe_451_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_483_io_input_valid = io_input_valid_483; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_483_io_iormac = io_iormac_483; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_484_clock = clock;
  assign bc_pe_484_reset = reset;
  assign bc_pe_484_io_ho_input = bc_pe_483_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_484_io_ve_input = bc_pe_452_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_484_io_input_valid = io_input_valid_484; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_484_io_iormac = io_iormac_484; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_485_clock = clock;
  assign bc_pe_485_reset = reset;
  assign bc_pe_485_io_ho_input = bc_pe_484_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_485_io_ve_input = bc_pe_453_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_485_io_input_valid = io_input_valid_485; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_485_io_iormac = io_iormac_485; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_486_clock = clock;
  assign bc_pe_486_reset = reset;
  assign bc_pe_486_io_ho_input = bc_pe_485_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_486_io_ve_input = bc_pe_454_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_486_io_input_valid = io_input_valid_486; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_486_io_iormac = io_iormac_486; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_487_clock = clock;
  assign bc_pe_487_reset = reset;
  assign bc_pe_487_io_ho_input = bc_pe_486_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_487_io_ve_input = bc_pe_455_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_487_io_input_valid = io_input_valid_487; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_487_io_iormac = io_iormac_487; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_488_clock = clock;
  assign bc_pe_488_reset = reset;
  assign bc_pe_488_io_ho_input = bc_pe_487_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_488_io_ve_input = bc_pe_456_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_488_io_input_valid = io_input_valid_488; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_488_io_iormac = io_iormac_488; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_489_clock = clock;
  assign bc_pe_489_reset = reset;
  assign bc_pe_489_io_ho_input = bc_pe_488_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_489_io_ve_input = bc_pe_457_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_489_io_input_valid = io_input_valid_489; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_489_io_iormac = io_iormac_489; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_490_clock = clock;
  assign bc_pe_490_reset = reset;
  assign bc_pe_490_io_ho_input = bc_pe_489_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_490_io_ve_input = bc_pe_458_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_490_io_input_valid = io_input_valid_490; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_490_io_iormac = io_iormac_490; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_491_clock = clock;
  assign bc_pe_491_reset = reset;
  assign bc_pe_491_io_ho_input = bc_pe_490_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_491_io_ve_input = bc_pe_459_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_491_io_input_valid = io_input_valid_491; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_491_io_iormac = io_iormac_491; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_492_clock = clock;
  assign bc_pe_492_reset = reset;
  assign bc_pe_492_io_ho_input = bc_pe_491_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_492_io_ve_input = bc_pe_460_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_492_io_input_valid = io_input_valid_492; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_492_io_iormac = io_iormac_492; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_493_clock = clock;
  assign bc_pe_493_reset = reset;
  assign bc_pe_493_io_ho_input = bc_pe_492_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_493_io_ve_input = bc_pe_461_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_493_io_input_valid = io_input_valid_493; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_493_io_iormac = io_iormac_493; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_494_clock = clock;
  assign bc_pe_494_reset = reset;
  assign bc_pe_494_io_ho_input = bc_pe_493_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_494_io_ve_input = bc_pe_462_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_494_io_input_valid = io_input_valid_494; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_494_io_iormac = io_iormac_494; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_495_clock = clock;
  assign bc_pe_495_reset = reset;
  assign bc_pe_495_io_ho_input = bc_pe_494_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_495_io_ve_input = bc_pe_463_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_495_io_input_valid = io_input_valid_495; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_495_io_iormac = io_iormac_495; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_496_clock = clock;
  assign bc_pe_496_reset = reset;
  assign bc_pe_496_io_ho_input = bc_pe_495_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_496_io_ve_input = bc_pe_464_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_496_io_input_valid = io_input_valid_496; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_496_io_iormac = io_iormac_496; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_497_clock = clock;
  assign bc_pe_497_reset = reset;
  assign bc_pe_497_io_ho_input = bc_pe_496_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_497_io_ve_input = bc_pe_465_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_497_io_input_valid = io_input_valid_497; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_497_io_iormac = io_iormac_497; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_498_clock = clock;
  assign bc_pe_498_reset = reset;
  assign bc_pe_498_io_ho_input = bc_pe_497_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_498_io_ve_input = bc_pe_466_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_498_io_input_valid = io_input_valid_498; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_498_io_iormac = io_iormac_498; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_499_clock = clock;
  assign bc_pe_499_reset = reset;
  assign bc_pe_499_io_ho_input = bc_pe_498_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_499_io_ve_input = bc_pe_467_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_499_io_input_valid = io_input_valid_499; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_499_io_iormac = io_iormac_499; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_500_clock = clock;
  assign bc_pe_500_reset = reset;
  assign bc_pe_500_io_ho_input = bc_pe_499_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_500_io_ve_input = bc_pe_468_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_500_io_input_valid = io_input_valid_500; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_500_io_iormac = io_iormac_500; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_501_clock = clock;
  assign bc_pe_501_reset = reset;
  assign bc_pe_501_io_ho_input = bc_pe_500_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_501_io_ve_input = bc_pe_469_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_501_io_input_valid = io_input_valid_501; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_501_io_iormac = io_iormac_501; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_502_clock = clock;
  assign bc_pe_502_reset = reset;
  assign bc_pe_502_io_ho_input = bc_pe_501_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_502_io_ve_input = bc_pe_470_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_502_io_input_valid = io_input_valid_502; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_502_io_iormac = io_iormac_502; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_503_clock = clock;
  assign bc_pe_503_reset = reset;
  assign bc_pe_503_io_ho_input = bc_pe_502_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_503_io_ve_input = bc_pe_471_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_503_io_input_valid = io_input_valid_503; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_503_io_iormac = io_iormac_503; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_504_clock = clock;
  assign bc_pe_504_reset = reset;
  assign bc_pe_504_io_ho_input = bc_pe_503_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_504_io_ve_input = bc_pe_472_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_504_io_input_valid = io_input_valid_504; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_504_io_iormac = io_iormac_504; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_505_clock = clock;
  assign bc_pe_505_reset = reset;
  assign bc_pe_505_io_ho_input = bc_pe_504_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_505_io_ve_input = bc_pe_473_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_505_io_input_valid = io_input_valid_505; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_505_io_iormac = io_iormac_505; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_506_clock = clock;
  assign bc_pe_506_reset = reset;
  assign bc_pe_506_io_ho_input = bc_pe_505_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_506_io_ve_input = bc_pe_474_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_506_io_input_valid = io_input_valid_506; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_506_io_iormac = io_iormac_506; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_507_clock = clock;
  assign bc_pe_507_reset = reset;
  assign bc_pe_507_io_ho_input = bc_pe_506_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_507_io_ve_input = bc_pe_475_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_507_io_input_valid = io_input_valid_507; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_507_io_iormac = io_iormac_507; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_508_clock = clock;
  assign bc_pe_508_reset = reset;
  assign bc_pe_508_io_ho_input = bc_pe_507_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_508_io_ve_input = bc_pe_476_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_508_io_input_valid = io_input_valid_508; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_508_io_iormac = io_iormac_508; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_509_clock = clock;
  assign bc_pe_509_reset = reset;
  assign bc_pe_509_io_ho_input = bc_pe_508_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_509_io_ve_input = bc_pe_477_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_509_io_input_valid = io_input_valid_509; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_509_io_iormac = io_iormac_509; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_510_clock = clock;
  assign bc_pe_510_reset = reset;
  assign bc_pe_510_io_ho_input = bc_pe_509_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_510_io_ve_input = bc_pe_478_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_510_io_input_valid = io_input_valid_510; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_510_io_iormac = io_iormac_510; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_511_clock = clock;
  assign bc_pe_511_reset = reset;
  assign bc_pe_511_io_ho_input = bc_pe_510_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_511_io_ve_input = bc_pe_479_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_511_io_input_valid = io_input_valid_511; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_511_io_iormac = io_iormac_511; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_512_clock = clock;
  assign bc_pe_512_reset = reset;
  assign bc_pe_512_io_ho_input = io_x_input_16; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_512_io_ve_input = bc_pe_480_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_512_io_input_valid = io_input_valid_512; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_512_io_iormac = io_iormac_512; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_513_clock = clock;
  assign bc_pe_513_reset = reset;
  assign bc_pe_513_io_ho_input = bc_pe_512_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_513_io_ve_input = bc_pe_481_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_513_io_input_valid = io_input_valid_513; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_513_io_iormac = io_iormac_513; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_514_clock = clock;
  assign bc_pe_514_reset = reset;
  assign bc_pe_514_io_ho_input = bc_pe_513_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_514_io_ve_input = bc_pe_482_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_514_io_input_valid = io_input_valid_514; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_514_io_iormac = io_iormac_514; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_515_clock = clock;
  assign bc_pe_515_reset = reset;
  assign bc_pe_515_io_ho_input = bc_pe_514_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_515_io_ve_input = bc_pe_483_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_515_io_input_valid = io_input_valid_515; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_515_io_iormac = io_iormac_515; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_516_clock = clock;
  assign bc_pe_516_reset = reset;
  assign bc_pe_516_io_ho_input = bc_pe_515_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_516_io_ve_input = bc_pe_484_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_516_io_input_valid = io_input_valid_516; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_516_io_iormac = io_iormac_516; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_517_clock = clock;
  assign bc_pe_517_reset = reset;
  assign bc_pe_517_io_ho_input = bc_pe_516_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_517_io_ve_input = bc_pe_485_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_517_io_input_valid = io_input_valid_517; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_517_io_iormac = io_iormac_517; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_518_clock = clock;
  assign bc_pe_518_reset = reset;
  assign bc_pe_518_io_ho_input = bc_pe_517_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_518_io_ve_input = bc_pe_486_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_518_io_input_valid = io_input_valid_518; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_518_io_iormac = io_iormac_518; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_519_clock = clock;
  assign bc_pe_519_reset = reset;
  assign bc_pe_519_io_ho_input = bc_pe_518_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_519_io_ve_input = bc_pe_487_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_519_io_input_valid = io_input_valid_519; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_519_io_iormac = io_iormac_519; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_520_clock = clock;
  assign bc_pe_520_reset = reset;
  assign bc_pe_520_io_ho_input = bc_pe_519_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_520_io_ve_input = bc_pe_488_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_520_io_input_valid = io_input_valid_520; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_520_io_iormac = io_iormac_520; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_521_clock = clock;
  assign bc_pe_521_reset = reset;
  assign bc_pe_521_io_ho_input = bc_pe_520_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_521_io_ve_input = bc_pe_489_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_521_io_input_valid = io_input_valid_521; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_521_io_iormac = io_iormac_521; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_522_clock = clock;
  assign bc_pe_522_reset = reset;
  assign bc_pe_522_io_ho_input = bc_pe_521_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_522_io_ve_input = bc_pe_490_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_522_io_input_valid = io_input_valid_522; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_522_io_iormac = io_iormac_522; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_523_clock = clock;
  assign bc_pe_523_reset = reset;
  assign bc_pe_523_io_ho_input = bc_pe_522_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_523_io_ve_input = bc_pe_491_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_523_io_input_valid = io_input_valid_523; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_523_io_iormac = io_iormac_523; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_524_clock = clock;
  assign bc_pe_524_reset = reset;
  assign bc_pe_524_io_ho_input = bc_pe_523_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_524_io_ve_input = bc_pe_492_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_524_io_input_valid = io_input_valid_524; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_524_io_iormac = io_iormac_524; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_525_clock = clock;
  assign bc_pe_525_reset = reset;
  assign bc_pe_525_io_ho_input = bc_pe_524_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_525_io_ve_input = bc_pe_493_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_525_io_input_valid = io_input_valid_525; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_525_io_iormac = io_iormac_525; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_526_clock = clock;
  assign bc_pe_526_reset = reset;
  assign bc_pe_526_io_ho_input = bc_pe_525_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_526_io_ve_input = bc_pe_494_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_526_io_input_valid = io_input_valid_526; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_526_io_iormac = io_iormac_526; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_527_clock = clock;
  assign bc_pe_527_reset = reset;
  assign bc_pe_527_io_ho_input = bc_pe_526_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_527_io_ve_input = bc_pe_495_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_527_io_input_valid = io_input_valid_527; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_527_io_iormac = io_iormac_527; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_528_clock = clock;
  assign bc_pe_528_reset = reset;
  assign bc_pe_528_io_ho_input = bc_pe_527_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_528_io_ve_input = bc_pe_496_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_528_io_input_valid = io_input_valid_528; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_528_io_iormac = io_iormac_528; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_529_clock = clock;
  assign bc_pe_529_reset = reset;
  assign bc_pe_529_io_ho_input = bc_pe_528_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_529_io_ve_input = bc_pe_497_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_529_io_input_valid = io_input_valid_529; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_529_io_iormac = io_iormac_529; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_530_clock = clock;
  assign bc_pe_530_reset = reset;
  assign bc_pe_530_io_ho_input = bc_pe_529_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_530_io_ve_input = bc_pe_498_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_530_io_input_valid = io_input_valid_530; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_530_io_iormac = io_iormac_530; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_531_clock = clock;
  assign bc_pe_531_reset = reset;
  assign bc_pe_531_io_ho_input = bc_pe_530_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_531_io_ve_input = bc_pe_499_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_531_io_input_valid = io_input_valid_531; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_531_io_iormac = io_iormac_531; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_532_clock = clock;
  assign bc_pe_532_reset = reset;
  assign bc_pe_532_io_ho_input = bc_pe_531_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_532_io_ve_input = bc_pe_500_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_532_io_input_valid = io_input_valid_532; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_532_io_iormac = io_iormac_532; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_533_clock = clock;
  assign bc_pe_533_reset = reset;
  assign bc_pe_533_io_ho_input = bc_pe_532_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_533_io_ve_input = bc_pe_501_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_533_io_input_valid = io_input_valid_533; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_533_io_iormac = io_iormac_533; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_534_clock = clock;
  assign bc_pe_534_reset = reset;
  assign bc_pe_534_io_ho_input = bc_pe_533_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_534_io_ve_input = bc_pe_502_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_534_io_input_valid = io_input_valid_534; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_534_io_iormac = io_iormac_534; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_535_clock = clock;
  assign bc_pe_535_reset = reset;
  assign bc_pe_535_io_ho_input = bc_pe_534_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_535_io_ve_input = bc_pe_503_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_535_io_input_valid = io_input_valid_535; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_535_io_iormac = io_iormac_535; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_536_clock = clock;
  assign bc_pe_536_reset = reset;
  assign bc_pe_536_io_ho_input = bc_pe_535_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_536_io_ve_input = bc_pe_504_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_536_io_input_valid = io_input_valid_536; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_536_io_iormac = io_iormac_536; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_537_clock = clock;
  assign bc_pe_537_reset = reset;
  assign bc_pe_537_io_ho_input = bc_pe_536_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_537_io_ve_input = bc_pe_505_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_537_io_input_valid = io_input_valid_537; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_537_io_iormac = io_iormac_537; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_538_clock = clock;
  assign bc_pe_538_reset = reset;
  assign bc_pe_538_io_ho_input = bc_pe_537_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_538_io_ve_input = bc_pe_506_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_538_io_input_valid = io_input_valid_538; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_538_io_iormac = io_iormac_538; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_539_clock = clock;
  assign bc_pe_539_reset = reset;
  assign bc_pe_539_io_ho_input = bc_pe_538_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_539_io_ve_input = bc_pe_507_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_539_io_input_valid = io_input_valid_539; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_539_io_iormac = io_iormac_539; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_540_clock = clock;
  assign bc_pe_540_reset = reset;
  assign bc_pe_540_io_ho_input = bc_pe_539_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_540_io_ve_input = bc_pe_508_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_540_io_input_valid = io_input_valid_540; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_540_io_iormac = io_iormac_540; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_541_clock = clock;
  assign bc_pe_541_reset = reset;
  assign bc_pe_541_io_ho_input = bc_pe_540_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_541_io_ve_input = bc_pe_509_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_541_io_input_valid = io_input_valid_541; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_541_io_iormac = io_iormac_541; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_542_clock = clock;
  assign bc_pe_542_reset = reset;
  assign bc_pe_542_io_ho_input = bc_pe_541_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_542_io_ve_input = bc_pe_510_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_542_io_input_valid = io_input_valid_542; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_542_io_iormac = io_iormac_542; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_543_clock = clock;
  assign bc_pe_543_reset = reset;
  assign bc_pe_543_io_ho_input = bc_pe_542_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_543_io_ve_input = bc_pe_511_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_543_io_input_valid = io_input_valid_543; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_543_io_iormac = io_iormac_543; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_544_clock = clock;
  assign bc_pe_544_reset = reset;
  assign bc_pe_544_io_ho_input = io_x_input_17; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_544_io_ve_input = bc_pe_512_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_544_io_input_valid = io_input_valid_544; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_544_io_iormac = io_iormac_544; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_545_clock = clock;
  assign bc_pe_545_reset = reset;
  assign bc_pe_545_io_ho_input = bc_pe_544_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_545_io_ve_input = bc_pe_513_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_545_io_input_valid = io_input_valid_545; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_545_io_iormac = io_iormac_545; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_546_clock = clock;
  assign bc_pe_546_reset = reset;
  assign bc_pe_546_io_ho_input = bc_pe_545_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_546_io_ve_input = bc_pe_514_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_546_io_input_valid = io_input_valid_546; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_546_io_iormac = io_iormac_546; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_547_clock = clock;
  assign bc_pe_547_reset = reset;
  assign bc_pe_547_io_ho_input = bc_pe_546_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_547_io_ve_input = bc_pe_515_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_547_io_input_valid = io_input_valid_547; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_547_io_iormac = io_iormac_547; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_548_clock = clock;
  assign bc_pe_548_reset = reset;
  assign bc_pe_548_io_ho_input = bc_pe_547_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_548_io_ve_input = bc_pe_516_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_548_io_input_valid = io_input_valid_548; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_548_io_iormac = io_iormac_548; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_549_clock = clock;
  assign bc_pe_549_reset = reset;
  assign bc_pe_549_io_ho_input = bc_pe_548_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_549_io_ve_input = bc_pe_517_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_549_io_input_valid = io_input_valid_549; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_549_io_iormac = io_iormac_549; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_550_clock = clock;
  assign bc_pe_550_reset = reset;
  assign bc_pe_550_io_ho_input = bc_pe_549_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_550_io_ve_input = bc_pe_518_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_550_io_input_valid = io_input_valid_550; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_550_io_iormac = io_iormac_550; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_551_clock = clock;
  assign bc_pe_551_reset = reset;
  assign bc_pe_551_io_ho_input = bc_pe_550_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_551_io_ve_input = bc_pe_519_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_551_io_input_valid = io_input_valid_551; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_551_io_iormac = io_iormac_551; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_552_clock = clock;
  assign bc_pe_552_reset = reset;
  assign bc_pe_552_io_ho_input = bc_pe_551_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_552_io_ve_input = bc_pe_520_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_552_io_input_valid = io_input_valid_552; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_552_io_iormac = io_iormac_552; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_553_clock = clock;
  assign bc_pe_553_reset = reset;
  assign bc_pe_553_io_ho_input = bc_pe_552_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_553_io_ve_input = bc_pe_521_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_553_io_input_valid = io_input_valid_553; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_553_io_iormac = io_iormac_553; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_554_clock = clock;
  assign bc_pe_554_reset = reset;
  assign bc_pe_554_io_ho_input = bc_pe_553_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_554_io_ve_input = bc_pe_522_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_554_io_input_valid = io_input_valid_554; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_554_io_iormac = io_iormac_554; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_555_clock = clock;
  assign bc_pe_555_reset = reset;
  assign bc_pe_555_io_ho_input = bc_pe_554_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_555_io_ve_input = bc_pe_523_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_555_io_input_valid = io_input_valid_555; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_555_io_iormac = io_iormac_555; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_556_clock = clock;
  assign bc_pe_556_reset = reset;
  assign bc_pe_556_io_ho_input = bc_pe_555_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_556_io_ve_input = bc_pe_524_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_556_io_input_valid = io_input_valid_556; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_556_io_iormac = io_iormac_556; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_557_clock = clock;
  assign bc_pe_557_reset = reset;
  assign bc_pe_557_io_ho_input = bc_pe_556_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_557_io_ve_input = bc_pe_525_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_557_io_input_valid = io_input_valid_557; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_557_io_iormac = io_iormac_557; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_558_clock = clock;
  assign bc_pe_558_reset = reset;
  assign bc_pe_558_io_ho_input = bc_pe_557_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_558_io_ve_input = bc_pe_526_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_558_io_input_valid = io_input_valid_558; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_558_io_iormac = io_iormac_558; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_559_clock = clock;
  assign bc_pe_559_reset = reset;
  assign bc_pe_559_io_ho_input = bc_pe_558_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_559_io_ve_input = bc_pe_527_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_559_io_input_valid = io_input_valid_559; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_559_io_iormac = io_iormac_559; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_560_clock = clock;
  assign bc_pe_560_reset = reset;
  assign bc_pe_560_io_ho_input = bc_pe_559_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_560_io_ve_input = bc_pe_528_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_560_io_input_valid = io_input_valid_560; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_560_io_iormac = io_iormac_560; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_561_clock = clock;
  assign bc_pe_561_reset = reset;
  assign bc_pe_561_io_ho_input = bc_pe_560_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_561_io_ve_input = bc_pe_529_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_561_io_input_valid = io_input_valid_561; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_561_io_iormac = io_iormac_561; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_562_clock = clock;
  assign bc_pe_562_reset = reset;
  assign bc_pe_562_io_ho_input = bc_pe_561_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_562_io_ve_input = bc_pe_530_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_562_io_input_valid = io_input_valid_562; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_562_io_iormac = io_iormac_562; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_563_clock = clock;
  assign bc_pe_563_reset = reset;
  assign bc_pe_563_io_ho_input = bc_pe_562_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_563_io_ve_input = bc_pe_531_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_563_io_input_valid = io_input_valid_563; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_563_io_iormac = io_iormac_563; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_564_clock = clock;
  assign bc_pe_564_reset = reset;
  assign bc_pe_564_io_ho_input = bc_pe_563_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_564_io_ve_input = bc_pe_532_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_564_io_input_valid = io_input_valid_564; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_564_io_iormac = io_iormac_564; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_565_clock = clock;
  assign bc_pe_565_reset = reset;
  assign bc_pe_565_io_ho_input = bc_pe_564_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_565_io_ve_input = bc_pe_533_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_565_io_input_valid = io_input_valid_565; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_565_io_iormac = io_iormac_565; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_566_clock = clock;
  assign bc_pe_566_reset = reset;
  assign bc_pe_566_io_ho_input = bc_pe_565_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_566_io_ve_input = bc_pe_534_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_566_io_input_valid = io_input_valid_566; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_566_io_iormac = io_iormac_566; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_567_clock = clock;
  assign bc_pe_567_reset = reset;
  assign bc_pe_567_io_ho_input = bc_pe_566_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_567_io_ve_input = bc_pe_535_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_567_io_input_valid = io_input_valid_567; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_567_io_iormac = io_iormac_567; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_568_clock = clock;
  assign bc_pe_568_reset = reset;
  assign bc_pe_568_io_ho_input = bc_pe_567_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_568_io_ve_input = bc_pe_536_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_568_io_input_valid = io_input_valid_568; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_568_io_iormac = io_iormac_568; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_569_clock = clock;
  assign bc_pe_569_reset = reset;
  assign bc_pe_569_io_ho_input = bc_pe_568_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_569_io_ve_input = bc_pe_537_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_569_io_input_valid = io_input_valid_569; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_569_io_iormac = io_iormac_569; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_570_clock = clock;
  assign bc_pe_570_reset = reset;
  assign bc_pe_570_io_ho_input = bc_pe_569_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_570_io_ve_input = bc_pe_538_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_570_io_input_valid = io_input_valid_570; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_570_io_iormac = io_iormac_570; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_571_clock = clock;
  assign bc_pe_571_reset = reset;
  assign bc_pe_571_io_ho_input = bc_pe_570_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_571_io_ve_input = bc_pe_539_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_571_io_input_valid = io_input_valid_571; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_571_io_iormac = io_iormac_571; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_572_clock = clock;
  assign bc_pe_572_reset = reset;
  assign bc_pe_572_io_ho_input = bc_pe_571_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_572_io_ve_input = bc_pe_540_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_572_io_input_valid = io_input_valid_572; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_572_io_iormac = io_iormac_572; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_573_clock = clock;
  assign bc_pe_573_reset = reset;
  assign bc_pe_573_io_ho_input = bc_pe_572_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_573_io_ve_input = bc_pe_541_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_573_io_input_valid = io_input_valid_573; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_573_io_iormac = io_iormac_573; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_574_clock = clock;
  assign bc_pe_574_reset = reset;
  assign bc_pe_574_io_ho_input = bc_pe_573_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_574_io_ve_input = bc_pe_542_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_574_io_input_valid = io_input_valid_574; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_574_io_iormac = io_iormac_574; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_575_clock = clock;
  assign bc_pe_575_reset = reset;
  assign bc_pe_575_io_ho_input = bc_pe_574_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_575_io_ve_input = bc_pe_543_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_575_io_input_valid = io_input_valid_575; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_575_io_iormac = io_iormac_575; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_576_clock = clock;
  assign bc_pe_576_reset = reset;
  assign bc_pe_576_io_ho_input = io_x_input_18; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_576_io_ve_input = bc_pe_544_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_576_io_input_valid = io_input_valid_576; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_576_io_iormac = io_iormac_576; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_577_clock = clock;
  assign bc_pe_577_reset = reset;
  assign bc_pe_577_io_ho_input = bc_pe_576_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_577_io_ve_input = bc_pe_545_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_577_io_input_valid = io_input_valid_577; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_577_io_iormac = io_iormac_577; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_578_clock = clock;
  assign bc_pe_578_reset = reset;
  assign bc_pe_578_io_ho_input = bc_pe_577_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_578_io_ve_input = bc_pe_546_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_578_io_input_valid = io_input_valid_578; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_578_io_iormac = io_iormac_578; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_579_clock = clock;
  assign bc_pe_579_reset = reset;
  assign bc_pe_579_io_ho_input = bc_pe_578_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_579_io_ve_input = bc_pe_547_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_579_io_input_valid = io_input_valid_579; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_579_io_iormac = io_iormac_579; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_580_clock = clock;
  assign bc_pe_580_reset = reset;
  assign bc_pe_580_io_ho_input = bc_pe_579_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_580_io_ve_input = bc_pe_548_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_580_io_input_valid = io_input_valid_580; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_580_io_iormac = io_iormac_580; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_581_clock = clock;
  assign bc_pe_581_reset = reset;
  assign bc_pe_581_io_ho_input = bc_pe_580_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_581_io_ve_input = bc_pe_549_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_581_io_input_valid = io_input_valid_581; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_581_io_iormac = io_iormac_581; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_582_clock = clock;
  assign bc_pe_582_reset = reset;
  assign bc_pe_582_io_ho_input = bc_pe_581_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_582_io_ve_input = bc_pe_550_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_582_io_input_valid = io_input_valid_582; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_582_io_iormac = io_iormac_582; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_583_clock = clock;
  assign bc_pe_583_reset = reset;
  assign bc_pe_583_io_ho_input = bc_pe_582_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_583_io_ve_input = bc_pe_551_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_583_io_input_valid = io_input_valid_583; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_583_io_iormac = io_iormac_583; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_584_clock = clock;
  assign bc_pe_584_reset = reset;
  assign bc_pe_584_io_ho_input = bc_pe_583_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_584_io_ve_input = bc_pe_552_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_584_io_input_valid = io_input_valid_584; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_584_io_iormac = io_iormac_584; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_585_clock = clock;
  assign bc_pe_585_reset = reset;
  assign bc_pe_585_io_ho_input = bc_pe_584_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_585_io_ve_input = bc_pe_553_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_585_io_input_valid = io_input_valid_585; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_585_io_iormac = io_iormac_585; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_586_clock = clock;
  assign bc_pe_586_reset = reset;
  assign bc_pe_586_io_ho_input = bc_pe_585_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_586_io_ve_input = bc_pe_554_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_586_io_input_valid = io_input_valid_586; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_586_io_iormac = io_iormac_586; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_587_clock = clock;
  assign bc_pe_587_reset = reset;
  assign bc_pe_587_io_ho_input = bc_pe_586_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_587_io_ve_input = bc_pe_555_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_587_io_input_valid = io_input_valid_587; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_587_io_iormac = io_iormac_587; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_588_clock = clock;
  assign bc_pe_588_reset = reset;
  assign bc_pe_588_io_ho_input = bc_pe_587_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_588_io_ve_input = bc_pe_556_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_588_io_input_valid = io_input_valid_588; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_588_io_iormac = io_iormac_588; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_589_clock = clock;
  assign bc_pe_589_reset = reset;
  assign bc_pe_589_io_ho_input = bc_pe_588_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_589_io_ve_input = bc_pe_557_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_589_io_input_valid = io_input_valid_589; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_589_io_iormac = io_iormac_589; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_590_clock = clock;
  assign bc_pe_590_reset = reset;
  assign bc_pe_590_io_ho_input = bc_pe_589_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_590_io_ve_input = bc_pe_558_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_590_io_input_valid = io_input_valid_590; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_590_io_iormac = io_iormac_590; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_591_clock = clock;
  assign bc_pe_591_reset = reset;
  assign bc_pe_591_io_ho_input = bc_pe_590_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_591_io_ve_input = bc_pe_559_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_591_io_input_valid = io_input_valid_591; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_591_io_iormac = io_iormac_591; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_592_clock = clock;
  assign bc_pe_592_reset = reset;
  assign bc_pe_592_io_ho_input = bc_pe_591_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_592_io_ve_input = bc_pe_560_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_592_io_input_valid = io_input_valid_592; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_592_io_iormac = io_iormac_592; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_593_clock = clock;
  assign bc_pe_593_reset = reset;
  assign bc_pe_593_io_ho_input = bc_pe_592_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_593_io_ve_input = bc_pe_561_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_593_io_input_valid = io_input_valid_593; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_593_io_iormac = io_iormac_593; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_594_clock = clock;
  assign bc_pe_594_reset = reset;
  assign bc_pe_594_io_ho_input = bc_pe_593_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_594_io_ve_input = bc_pe_562_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_594_io_input_valid = io_input_valid_594; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_594_io_iormac = io_iormac_594; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_595_clock = clock;
  assign bc_pe_595_reset = reset;
  assign bc_pe_595_io_ho_input = bc_pe_594_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_595_io_ve_input = bc_pe_563_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_595_io_input_valid = io_input_valid_595; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_595_io_iormac = io_iormac_595; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_596_clock = clock;
  assign bc_pe_596_reset = reset;
  assign bc_pe_596_io_ho_input = bc_pe_595_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_596_io_ve_input = bc_pe_564_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_596_io_input_valid = io_input_valid_596; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_596_io_iormac = io_iormac_596; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_597_clock = clock;
  assign bc_pe_597_reset = reset;
  assign bc_pe_597_io_ho_input = bc_pe_596_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_597_io_ve_input = bc_pe_565_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_597_io_input_valid = io_input_valid_597; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_597_io_iormac = io_iormac_597; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_598_clock = clock;
  assign bc_pe_598_reset = reset;
  assign bc_pe_598_io_ho_input = bc_pe_597_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_598_io_ve_input = bc_pe_566_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_598_io_input_valid = io_input_valid_598; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_598_io_iormac = io_iormac_598; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_599_clock = clock;
  assign bc_pe_599_reset = reset;
  assign bc_pe_599_io_ho_input = bc_pe_598_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_599_io_ve_input = bc_pe_567_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_599_io_input_valid = io_input_valid_599; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_599_io_iormac = io_iormac_599; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_600_clock = clock;
  assign bc_pe_600_reset = reset;
  assign bc_pe_600_io_ho_input = bc_pe_599_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_600_io_ve_input = bc_pe_568_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_600_io_input_valid = io_input_valid_600; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_600_io_iormac = io_iormac_600; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_601_clock = clock;
  assign bc_pe_601_reset = reset;
  assign bc_pe_601_io_ho_input = bc_pe_600_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_601_io_ve_input = bc_pe_569_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_601_io_input_valid = io_input_valid_601; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_601_io_iormac = io_iormac_601; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_602_clock = clock;
  assign bc_pe_602_reset = reset;
  assign bc_pe_602_io_ho_input = bc_pe_601_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_602_io_ve_input = bc_pe_570_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_602_io_input_valid = io_input_valid_602; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_602_io_iormac = io_iormac_602; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_603_clock = clock;
  assign bc_pe_603_reset = reset;
  assign bc_pe_603_io_ho_input = bc_pe_602_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_603_io_ve_input = bc_pe_571_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_603_io_input_valid = io_input_valid_603; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_603_io_iormac = io_iormac_603; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_604_clock = clock;
  assign bc_pe_604_reset = reset;
  assign bc_pe_604_io_ho_input = bc_pe_603_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_604_io_ve_input = bc_pe_572_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_604_io_input_valid = io_input_valid_604; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_604_io_iormac = io_iormac_604; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_605_clock = clock;
  assign bc_pe_605_reset = reset;
  assign bc_pe_605_io_ho_input = bc_pe_604_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_605_io_ve_input = bc_pe_573_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_605_io_input_valid = io_input_valid_605; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_605_io_iormac = io_iormac_605; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_606_clock = clock;
  assign bc_pe_606_reset = reset;
  assign bc_pe_606_io_ho_input = bc_pe_605_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_606_io_ve_input = bc_pe_574_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_606_io_input_valid = io_input_valid_606; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_606_io_iormac = io_iormac_606; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_607_clock = clock;
  assign bc_pe_607_reset = reset;
  assign bc_pe_607_io_ho_input = bc_pe_606_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_607_io_ve_input = bc_pe_575_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_607_io_input_valid = io_input_valid_607; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_607_io_iormac = io_iormac_607; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_608_clock = clock;
  assign bc_pe_608_reset = reset;
  assign bc_pe_608_io_ho_input = io_x_input_19; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_608_io_ve_input = bc_pe_576_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_608_io_input_valid = io_input_valid_608; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_608_io_iormac = io_iormac_608; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_609_clock = clock;
  assign bc_pe_609_reset = reset;
  assign bc_pe_609_io_ho_input = bc_pe_608_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_609_io_ve_input = bc_pe_577_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_609_io_input_valid = io_input_valid_609; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_609_io_iormac = io_iormac_609; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_610_clock = clock;
  assign bc_pe_610_reset = reset;
  assign bc_pe_610_io_ho_input = bc_pe_609_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_610_io_ve_input = bc_pe_578_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_610_io_input_valid = io_input_valid_610; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_610_io_iormac = io_iormac_610; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_611_clock = clock;
  assign bc_pe_611_reset = reset;
  assign bc_pe_611_io_ho_input = bc_pe_610_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_611_io_ve_input = bc_pe_579_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_611_io_input_valid = io_input_valid_611; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_611_io_iormac = io_iormac_611; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_612_clock = clock;
  assign bc_pe_612_reset = reset;
  assign bc_pe_612_io_ho_input = bc_pe_611_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_612_io_ve_input = bc_pe_580_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_612_io_input_valid = io_input_valid_612; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_612_io_iormac = io_iormac_612; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_613_clock = clock;
  assign bc_pe_613_reset = reset;
  assign bc_pe_613_io_ho_input = bc_pe_612_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_613_io_ve_input = bc_pe_581_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_613_io_input_valid = io_input_valid_613; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_613_io_iormac = io_iormac_613; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_614_clock = clock;
  assign bc_pe_614_reset = reset;
  assign bc_pe_614_io_ho_input = bc_pe_613_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_614_io_ve_input = bc_pe_582_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_614_io_input_valid = io_input_valid_614; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_614_io_iormac = io_iormac_614; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_615_clock = clock;
  assign bc_pe_615_reset = reset;
  assign bc_pe_615_io_ho_input = bc_pe_614_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_615_io_ve_input = bc_pe_583_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_615_io_input_valid = io_input_valid_615; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_615_io_iormac = io_iormac_615; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_616_clock = clock;
  assign bc_pe_616_reset = reset;
  assign bc_pe_616_io_ho_input = bc_pe_615_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_616_io_ve_input = bc_pe_584_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_616_io_input_valid = io_input_valid_616; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_616_io_iormac = io_iormac_616; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_617_clock = clock;
  assign bc_pe_617_reset = reset;
  assign bc_pe_617_io_ho_input = bc_pe_616_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_617_io_ve_input = bc_pe_585_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_617_io_input_valid = io_input_valid_617; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_617_io_iormac = io_iormac_617; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_618_clock = clock;
  assign bc_pe_618_reset = reset;
  assign bc_pe_618_io_ho_input = bc_pe_617_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_618_io_ve_input = bc_pe_586_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_618_io_input_valid = io_input_valid_618; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_618_io_iormac = io_iormac_618; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_619_clock = clock;
  assign bc_pe_619_reset = reset;
  assign bc_pe_619_io_ho_input = bc_pe_618_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_619_io_ve_input = bc_pe_587_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_619_io_input_valid = io_input_valid_619; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_619_io_iormac = io_iormac_619; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_620_clock = clock;
  assign bc_pe_620_reset = reset;
  assign bc_pe_620_io_ho_input = bc_pe_619_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_620_io_ve_input = bc_pe_588_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_620_io_input_valid = io_input_valid_620; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_620_io_iormac = io_iormac_620; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_621_clock = clock;
  assign bc_pe_621_reset = reset;
  assign bc_pe_621_io_ho_input = bc_pe_620_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_621_io_ve_input = bc_pe_589_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_621_io_input_valid = io_input_valid_621; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_621_io_iormac = io_iormac_621; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_622_clock = clock;
  assign bc_pe_622_reset = reset;
  assign bc_pe_622_io_ho_input = bc_pe_621_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_622_io_ve_input = bc_pe_590_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_622_io_input_valid = io_input_valid_622; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_622_io_iormac = io_iormac_622; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_623_clock = clock;
  assign bc_pe_623_reset = reset;
  assign bc_pe_623_io_ho_input = bc_pe_622_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_623_io_ve_input = bc_pe_591_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_623_io_input_valid = io_input_valid_623; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_623_io_iormac = io_iormac_623; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_624_clock = clock;
  assign bc_pe_624_reset = reset;
  assign bc_pe_624_io_ho_input = bc_pe_623_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_624_io_ve_input = bc_pe_592_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_624_io_input_valid = io_input_valid_624; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_624_io_iormac = io_iormac_624; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_625_clock = clock;
  assign bc_pe_625_reset = reset;
  assign bc_pe_625_io_ho_input = bc_pe_624_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_625_io_ve_input = bc_pe_593_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_625_io_input_valid = io_input_valid_625; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_625_io_iormac = io_iormac_625; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_626_clock = clock;
  assign bc_pe_626_reset = reset;
  assign bc_pe_626_io_ho_input = bc_pe_625_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_626_io_ve_input = bc_pe_594_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_626_io_input_valid = io_input_valid_626; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_626_io_iormac = io_iormac_626; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_627_clock = clock;
  assign bc_pe_627_reset = reset;
  assign bc_pe_627_io_ho_input = bc_pe_626_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_627_io_ve_input = bc_pe_595_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_627_io_input_valid = io_input_valid_627; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_627_io_iormac = io_iormac_627; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_628_clock = clock;
  assign bc_pe_628_reset = reset;
  assign bc_pe_628_io_ho_input = bc_pe_627_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_628_io_ve_input = bc_pe_596_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_628_io_input_valid = io_input_valid_628; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_628_io_iormac = io_iormac_628; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_629_clock = clock;
  assign bc_pe_629_reset = reset;
  assign bc_pe_629_io_ho_input = bc_pe_628_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_629_io_ve_input = bc_pe_597_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_629_io_input_valid = io_input_valid_629; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_629_io_iormac = io_iormac_629; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_630_clock = clock;
  assign bc_pe_630_reset = reset;
  assign bc_pe_630_io_ho_input = bc_pe_629_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_630_io_ve_input = bc_pe_598_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_630_io_input_valid = io_input_valid_630; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_630_io_iormac = io_iormac_630; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_631_clock = clock;
  assign bc_pe_631_reset = reset;
  assign bc_pe_631_io_ho_input = bc_pe_630_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_631_io_ve_input = bc_pe_599_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_631_io_input_valid = io_input_valid_631; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_631_io_iormac = io_iormac_631; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_632_clock = clock;
  assign bc_pe_632_reset = reset;
  assign bc_pe_632_io_ho_input = bc_pe_631_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_632_io_ve_input = bc_pe_600_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_632_io_input_valid = io_input_valid_632; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_632_io_iormac = io_iormac_632; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_633_clock = clock;
  assign bc_pe_633_reset = reset;
  assign bc_pe_633_io_ho_input = bc_pe_632_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_633_io_ve_input = bc_pe_601_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_633_io_input_valid = io_input_valid_633; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_633_io_iormac = io_iormac_633; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_634_clock = clock;
  assign bc_pe_634_reset = reset;
  assign bc_pe_634_io_ho_input = bc_pe_633_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_634_io_ve_input = bc_pe_602_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_634_io_input_valid = io_input_valid_634; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_634_io_iormac = io_iormac_634; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_635_clock = clock;
  assign bc_pe_635_reset = reset;
  assign bc_pe_635_io_ho_input = bc_pe_634_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_635_io_ve_input = bc_pe_603_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_635_io_input_valid = io_input_valid_635; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_635_io_iormac = io_iormac_635; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_636_clock = clock;
  assign bc_pe_636_reset = reset;
  assign bc_pe_636_io_ho_input = bc_pe_635_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_636_io_ve_input = bc_pe_604_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_636_io_input_valid = io_input_valid_636; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_636_io_iormac = io_iormac_636; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_637_clock = clock;
  assign bc_pe_637_reset = reset;
  assign bc_pe_637_io_ho_input = bc_pe_636_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_637_io_ve_input = bc_pe_605_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_637_io_input_valid = io_input_valid_637; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_637_io_iormac = io_iormac_637; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_638_clock = clock;
  assign bc_pe_638_reset = reset;
  assign bc_pe_638_io_ho_input = bc_pe_637_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_638_io_ve_input = bc_pe_606_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_638_io_input_valid = io_input_valid_638; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_638_io_iormac = io_iormac_638; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_639_clock = clock;
  assign bc_pe_639_reset = reset;
  assign bc_pe_639_io_ho_input = bc_pe_638_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_639_io_ve_input = bc_pe_607_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_639_io_input_valid = io_input_valid_639; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_639_io_iormac = io_iormac_639; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_640_clock = clock;
  assign bc_pe_640_reset = reset;
  assign bc_pe_640_io_ho_input = io_x_input_20; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_640_io_ve_input = bc_pe_608_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_640_io_input_valid = io_input_valid_640; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_640_io_iormac = io_iormac_640; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_641_clock = clock;
  assign bc_pe_641_reset = reset;
  assign bc_pe_641_io_ho_input = bc_pe_640_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_641_io_ve_input = bc_pe_609_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_641_io_input_valid = io_input_valid_641; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_641_io_iormac = io_iormac_641; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_642_clock = clock;
  assign bc_pe_642_reset = reset;
  assign bc_pe_642_io_ho_input = bc_pe_641_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_642_io_ve_input = bc_pe_610_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_642_io_input_valid = io_input_valid_642; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_642_io_iormac = io_iormac_642; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_643_clock = clock;
  assign bc_pe_643_reset = reset;
  assign bc_pe_643_io_ho_input = bc_pe_642_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_643_io_ve_input = bc_pe_611_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_643_io_input_valid = io_input_valid_643; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_643_io_iormac = io_iormac_643; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_644_clock = clock;
  assign bc_pe_644_reset = reset;
  assign bc_pe_644_io_ho_input = bc_pe_643_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_644_io_ve_input = bc_pe_612_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_644_io_input_valid = io_input_valid_644; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_644_io_iormac = io_iormac_644; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_645_clock = clock;
  assign bc_pe_645_reset = reset;
  assign bc_pe_645_io_ho_input = bc_pe_644_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_645_io_ve_input = bc_pe_613_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_645_io_input_valid = io_input_valid_645; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_645_io_iormac = io_iormac_645; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_646_clock = clock;
  assign bc_pe_646_reset = reset;
  assign bc_pe_646_io_ho_input = bc_pe_645_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_646_io_ve_input = bc_pe_614_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_646_io_input_valid = io_input_valid_646; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_646_io_iormac = io_iormac_646; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_647_clock = clock;
  assign bc_pe_647_reset = reset;
  assign bc_pe_647_io_ho_input = bc_pe_646_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_647_io_ve_input = bc_pe_615_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_647_io_input_valid = io_input_valid_647; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_647_io_iormac = io_iormac_647; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_648_clock = clock;
  assign bc_pe_648_reset = reset;
  assign bc_pe_648_io_ho_input = bc_pe_647_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_648_io_ve_input = bc_pe_616_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_648_io_input_valid = io_input_valid_648; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_648_io_iormac = io_iormac_648; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_649_clock = clock;
  assign bc_pe_649_reset = reset;
  assign bc_pe_649_io_ho_input = bc_pe_648_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_649_io_ve_input = bc_pe_617_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_649_io_input_valid = io_input_valid_649; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_649_io_iormac = io_iormac_649; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_650_clock = clock;
  assign bc_pe_650_reset = reset;
  assign bc_pe_650_io_ho_input = bc_pe_649_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_650_io_ve_input = bc_pe_618_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_650_io_input_valid = io_input_valid_650; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_650_io_iormac = io_iormac_650; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_651_clock = clock;
  assign bc_pe_651_reset = reset;
  assign bc_pe_651_io_ho_input = bc_pe_650_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_651_io_ve_input = bc_pe_619_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_651_io_input_valid = io_input_valid_651; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_651_io_iormac = io_iormac_651; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_652_clock = clock;
  assign bc_pe_652_reset = reset;
  assign bc_pe_652_io_ho_input = bc_pe_651_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_652_io_ve_input = bc_pe_620_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_652_io_input_valid = io_input_valid_652; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_652_io_iormac = io_iormac_652; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_653_clock = clock;
  assign bc_pe_653_reset = reset;
  assign bc_pe_653_io_ho_input = bc_pe_652_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_653_io_ve_input = bc_pe_621_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_653_io_input_valid = io_input_valid_653; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_653_io_iormac = io_iormac_653; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_654_clock = clock;
  assign bc_pe_654_reset = reset;
  assign bc_pe_654_io_ho_input = bc_pe_653_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_654_io_ve_input = bc_pe_622_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_654_io_input_valid = io_input_valid_654; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_654_io_iormac = io_iormac_654; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_655_clock = clock;
  assign bc_pe_655_reset = reset;
  assign bc_pe_655_io_ho_input = bc_pe_654_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_655_io_ve_input = bc_pe_623_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_655_io_input_valid = io_input_valid_655; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_655_io_iormac = io_iormac_655; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_656_clock = clock;
  assign bc_pe_656_reset = reset;
  assign bc_pe_656_io_ho_input = bc_pe_655_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_656_io_ve_input = bc_pe_624_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_656_io_input_valid = io_input_valid_656; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_656_io_iormac = io_iormac_656; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_657_clock = clock;
  assign bc_pe_657_reset = reset;
  assign bc_pe_657_io_ho_input = bc_pe_656_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_657_io_ve_input = bc_pe_625_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_657_io_input_valid = io_input_valid_657; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_657_io_iormac = io_iormac_657; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_658_clock = clock;
  assign bc_pe_658_reset = reset;
  assign bc_pe_658_io_ho_input = bc_pe_657_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_658_io_ve_input = bc_pe_626_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_658_io_input_valid = io_input_valid_658; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_658_io_iormac = io_iormac_658; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_659_clock = clock;
  assign bc_pe_659_reset = reset;
  assign bc_pe_659_io_ho_input = bc_pe_658_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_659_io_ve_input = bc_pe_627_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_659_io_input_valid = io_input_valid_659; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_659_io_iormac = io_iormac_659; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_660_clock = clock;
  assign bc_pe_660_reset = reset;
  assign bc_pe_660_io_ho_input = bc_pe_659_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_660_io_ve_input = bc_pe_628_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_660_io_input_valid = io_input_valid_660; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_660_io_iormac = io_iormac_660; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_661_clock = clock;
  assign bc_pe_661_reset = reset;
  assign bc_pe_661_io_ho_input = bc_pe_660_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_661_io_ve_input = bc_pe_629_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_661_io_input_valid = io_input_valid_661; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_661_io_iormac = io_iormac_661; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_662_clock = clock;
  assign bc_pe_662_reset = reset;
  assign bc_pe_662_io_ho_input = bc_pe_661_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_662_io_ve_input = bc_pe_630_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_662_io_input_valid = io_input_valid_662; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_662_io_iormac = io_iormac_662; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_663_clock = clock;
  assign bc_pe_663_reset = reset;
  assign bc_pe_663_io_ho_input = bc_pe_662_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_663_io_ve_input = bc_pe_631_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_663_io_input_valid = io_input_valid_663; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_663_io_iormac = io_iormac_663; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_664_clock = clock;
  assign bc_pe_664_reset = reset;
  assign bc_pe_664_io_ho_input = bc_pe_663_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_664_io_ve_input = bc_pe_632_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_664_io_input_valid = io_input_valid_664; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_664_io_iormac = io_iormac_664; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_665_clock = clock;
  assign bc_pe_665_reset = reset;
  assign bc_pe_665_io_ho_input = bc_pe_664_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_665_io_ve_input = bc_pe_633_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_665_io_input_valid = io_input_valid_665; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_665_io_iormac = io_iormac_665; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_666_clock = clock;
  assign bc_pe_666_reset = reset;
  assign bc_pe_666_io_ho_input = bc_pe_665_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_666_io_ve_input = bc_pe_634_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_666_io_input_valid = io_input_valid_666; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_666_io_iormac = io_iormac_666; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_667_clock = clock;
  assign bc_pe_667_reset = reset;
  assign bc_pe_667_io_ho_input = bc_pe_666_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_667_io_ve_input = bc_pe_635_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_667_io_input_valid = io_input_valid_667; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_667_io_iormac = io_iormac_667; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_668_clock = clock;
  assign bc_pe_668_reset = reset;
  assign bc_pe_668_io_ho_input = bc_pe_667_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_668_io_ve_input = bc_pe_636_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_668_io_input_valid = io_input_valid_668; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_668_io_iormac = io_iormac_668; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_669_clock = clock;
  assign bc_pe_669_reset = reset;
  assign bc_pe_669_io_ho_input = bc_pe_668_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_669_io_ve_input = bc_pe_637_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_669_io_input_valid = io_input_valid_669; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_669_io_iormac = io_iormac_669; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_670_clock = clock;
  assign bc_pe_670_reset = reset;
  assign bc_pe_670_io_ho_input = bc_pe_669_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_670_io_ve_input = bc_pe_638_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_670_io_input_valid = io_input_valid_670; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_670_io_iormac = io_iormac_670; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_671_clock = clock;
  assign bc_pe_671_reset = reset;
  assign bc_pe_671_io_ho_input = bc_pe_670_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_671_io_ve_input = bc_pe_639_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_671_io_input_valid = io_input_valid_671; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_671_io_iormac = io_iormac_671; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_672_clock = clock;
  assign bc_pe_672_reset = reset;
  assign bc_pe_672_io_ho_input = io_x_input_21; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_672_io_ve_input = bc_pe_640_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_672_io_input_valid = io_input_valid_672; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_672_io_iormac = io_iormac_672; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_673_clock = clock;
  assign bc_pe_673_reset = reset;
  assign bc_pe_673_io_ho_input = bc_pe_672_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_673_io_ve_input = bc_pe_641_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_673_io_input_valid = io_input_valid_673; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_673_io_iormac = io_iormac_673; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_674_clock = clock;
  assign bc_pe_674_reset = reset;
  assign bc_pe_674_io_ho_input = bc_pe_673_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_674_io_ve_input = bc_pe_642_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_674_io_input_valid = io_input_valid_674; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_674_io_iormac = io_iormac_674; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_675_clock = clock;
  assign bc_pe_675_reset = reset;
  assign bc_pe_675_io_ho_input = bc_pe_674_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_675_io_ve_input = bc_pe_643_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_675_io_input_valid = io_input_valid_675; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_675_io_iormac = io_iormac_675; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_676_clock = clock;
  assign bc_pe_676_reset = reset;
  assign bc_pe_676_io_ho_input = bc_pe_675_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_676_io_ve_input = bc_pe_644_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_676_io_input_valid = io_input_valid_676; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_676_io_iormac = io_iormac_676; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_677_clock = clock;
  assign bc_pe_677_reset = reset;
  assign bc_pe_677_io_ho_input = bc_pe_676_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_677_io_ve_input = bc_pe_645_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_677_io_input_valid = io_input_valid_677; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_677_io_iormac = io_iormac_677; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_678_clock = clock;
  assign bc_pe_678_reset = reset;
  assign bc_pe_678_io_ho_input = bc_pe_677_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_678_io_ve_input = bc_pe_646_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_678_io_input_valid = io_input_valid_678; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_678_io_iormac = io_iormac_678; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_679_clock = clock;
  assign bc_pe_679_reset = reset;
  assign bc_pe_679_io_ho_input = bc_pe_678_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_679_io_ve_input = bc_pe_647_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_679_io_input_valid = io_input_valid_679; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_679_io_iormac = io_iormac_679; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_680_clock = clock;
  assign bc_pe_680_reset = reset;
  assign bc_pe_680_io_ho_input = bc_pe_679_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_680_io_ve_input = bc_pe_648_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_680_io_input_valid = io_input_valid_680; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_680_io_iormac = io_iormac_680; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_681_clock = clock;
  assign bc_pe_681_reset = reset;
  assign bc_pe_681_io_ho_input = bc_pe_680_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_681_io_ve_input = bc_pe_649_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_681_io_input_valid = io_input_valid_681; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_681_io_iormac = io_iormac_681; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_682_clock = clock;
  assign bc_pe_682_reset = reset;
  assign bc_pe_682_io_ho_input = bc_pe_681_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_682_io_ve_input = bc_pe_650_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_682_io_input_valid = io_input_valid_682; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_682_io_iormac = io_iormac_682; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_683_clock = clock;
  assign bc_pe_683_reset = reset;
  assign bc_pe_683_io_ho_input = bc_pe_682_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_683_io_ve_input = bc_pe_651_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_683_io_input_valid = io_input_valid_683; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_683_io_iormac = io_iormac_683; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_684_clock = clock;
  assign bc_pe_684_reset = reset;
  assign bc_pe_684_io_ho_input = bc_pe_683_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_684_io_ve_input = bc_pe_652_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_684_io_input_valid = io_input_valid_684; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_684_io_iormac = io_iormac_684; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_685_clock = clock;
  assign bc_pe_685_reset = reset;
  assign bc_pe_685_io_ho_input = bc_pe_684_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_685_io_ve_input = bc_pe_653_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_685_io_input_valid = io_input_valid_685; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_685_io_iormac = io_iormac_685; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_686_clock = clock;
  assign bc_pe_686_reset = reset;
  assign bc_pe_686_io_ho_input = bc_pe_685_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_686_io_ve_input = bc_pe_654_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_686_io_input_valid = io_input_valid_686; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_686_io_iormac = io_iormac_686; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_687_clock = clock;
  assign bc_pe_687_reset = reset;
  assign bc_pe_687_io_ho_input = bc_pe_686_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_687_io_ve_input = bc_pe_655_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_687_io_input_valid = io_input_valid_687; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_687_io_iormac = io_iormac_687; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_688_clock = clock;
  assign bc_pe_688_reset = reset;
  assign bc_pe_688_io_ho_input = bc_pe_687_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_688_io_ve_input = bc_pe_656_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_688_io_input_valid = io_input_valid_688; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_688_io_iormac = io_iormac_688; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_689_clock = clock;
  assign bc_pe_689_reset = reset;
  assign bc_pe_689_io_ho_input = bc_pe_688_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_689_io_ve_input = bc_pe_657_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_689_io_input_valid = io_input_valid_689; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_689_io_iormac = io_iormac_689; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_690_clock = clock;
  assign bc_pe_690_reset = reset;
  assign bc_pe_690_io_ho_input = bc_pe_689_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_690_io_ve_input = bc_pe_658_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_690_io_input_valid = io_input_valid_690; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_690_io_iormac = io_iormac_690; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_691_clock = clock;
  assign bc_pe_691_reset = reset;
  assign bc_pe_691_io_ho_input = bc_pe_690_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_691_io_ve_input = bc_pe_659_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_691_io_input_valid = io_input_valid_691; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_691_io_iormac = io_iormac_691; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_692_clock = clock;
  assign bc_pe_692_reset = reset;
  assign bc_pe_692_io_ho_input = bc_pe_691_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_692_io_ve_input = bc_pe_660_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_692_io_input_valid = io_input_valid_692; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_692_io_iormac = io_iormac_692; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_693_clock = clock;
  assign bc_pe_693_reset = reset;
  assign bc_pe_693_io_ho_input = bc_pe_692_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_693_io_ve_input = bc_pe_661_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_693_io_input_valid = io_input_valid_693; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_693_io_iormac = io_iormac_693; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_694_clock = clock;
  assign bc_pe_694_reset = reset;
  assign bc_pe_694_io_ho_input = bc_pe_693_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_694_io_ve_input = bc_pe_662_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_694_io_input_valid = io_input_valid_694; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_694_io_iormac = io_iormac_694; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_695_clock = clock;
  assign bc_pe_695_reset = reset;
  assign bc_pe_695_io_ho_input = bc_pe_694_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_695_io_ve_input = bc_pe_663_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_695_io_input_valid = io_input_valid_695; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_695_io_iormac = io_iormac_695; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_696_clock = clock;
  assign bc_pe_696_reset = reset;
  assign bc_pe_696_io_ho_input = bc_pe_695_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_696_io_ve_input = bc_pe_664_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_696_io_input_valid = io_input_valid_696; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_696_io_iormac = io_iormac_696; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_697_clock = clock;
  assign bc_pe_697_reset = reset;
  assign bc_pe_697_io_ho_input = bc_pe_696_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_697_io_ve_input = bc_pe_665_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_697_io_input_valid = io_input_valid_697; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_697_io_iormac = io_iormac_697; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_698_clock = clock;
  assign bc_pe_698_reset = reset;
  assign bc_pe_698_io_ho_input = bc_pe_697_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_698_io_ve_input = bc_pe_666_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_698_io_input_valid = io_input_valid_698; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_698_io_iormac = io_iormac_698; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_699_clock = clock;
  assign bc_pe_699_reset = reset;
  assign bc_pe_699_io_ho_input = bc_pe_698_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_699_io_ve_input = bc_pe_667_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_699_io_input_valid = io_input_valid_699; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_699_io_iormac = io_iormac_699; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_700_clock = clock;
  assign bc_pe_700_reset = reset;
  assign bc_pe_700_io_ho_input = bc_pe_699_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_700_io_ve_input = bc_pe_668_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_700_io_input_valid = io_input_valid_700; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_700_io_iormac = io_iormac_700; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_701_clock = clock;
  assign bc_pe_701_reset = reset;
  assign bc_pe_701_io_ho_input = bc_pe_700_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_701_io_ve_input = bc_pe_669_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_701_io_input_valid = io_input_valid_701; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_701_io_iormac = io_iormac_701; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_702_clock = clock;
  assign bc_pe_702_reset = reset;
  assign bc_pe_702_io_ho_input = bc_pe_701_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_702_io_ve_input = bc_pe_670_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_702_io_input_valid = io_input_valid_702; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_702_io_iormac = io_iormac_702; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_703_clock = clock;
  assign bc_pe_703_reset = reset;
  assign bc_pe_703_io_ho_input = bc_pe_702_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_703_io_ve_input = bc_pe_671_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_703_io_input_valid = io_input_valid_703; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_703_io_iormac = io_iormac_703; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_704_clock = clock;
  assign bc_pe_704_reset = reset;
  assign bc_pe_704_io_ho_input = io_x_input_22; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_704_io_ve_input = bc_pe_672_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_704_io_input_valid = io_input_valid_704; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_704_io_iormac = io_iormac_704; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_705_clock = clock;
  assign bc_pe_705_reset = reset;
  assign bc_pe_705_io_ho_input = bc_pe_704_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_705_io_ve_input = bc_pe_673_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_705_io_input_valid = io_input_valid_705; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_705_io_iormac = io_iormac_705; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_706_clock = clock;
  assign bc_pe_706_reset = reset;
  assign bc_pe_706_io_ho_input = bc_pe_705_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_706_io_ve_input = bc_pe_674_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_706_io_input_valid = io_input_valid_706; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_706_io_iormac = io_iormac_706; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_707_clock = clock;
  assign bc_pe_707_reset = reset;
  assign bc_pe_707_io_ho_input = bc_pe_706_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_707_io_ve_input = bc_pe_675_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_707_io_input_valid = io_input_valid_707; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_707_io_iormac = io_iormac_707; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_708_clock = clock;
  assign bc_pe_708_reset = reset;
  assign bc_pe_708_io_ho_input = bc_pe_707_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_708_io_ve_input = bc_pe_676_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_708_io_input_valid = io_input_valid_708; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_708_io_iormac = io_iormac_708; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_709_clock = clock;
  assign bc_pe_709_reset = reset;
  assign bc_pe_709_io_ho_input = bc_pe_708_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_709_io_ve_input = bc_pe_677_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_709_io_input_valid = io_input_valid_709; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_709_io_iormac = io_iormac_709; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_710_clock = clock;
  assign bc_pe_710_reset = reset;
  assign bc_pe_710_io_ho_input = bc_pe_709_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_710_io_ve_input = bc_pe_678_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_710_io_input_valid = io_input_valid_710; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_710_io_iormac = io_iormac_710; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_711_clock = clock;
  assign bc_pe_711_reset = reset;
  assign bc_pe_711_io_ho_input = bc_pe_710_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_711_io_ve_input = bc_pe_679_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_711_io_input_valid = io_input_valid_711; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_711_io_iormac = io_iormac_711; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_712_clock = clock;
  assign bc_pe_712_reset = reset;
  assign bc_pe_712_io_ho_input = bc_pe_711_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_712_io_ve_input = bc_pe_680_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_712_io_input_valid = io_input_valid_712; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_712_io_iormac = io_iormac_712; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_713_clock = clock;
  assign bc_pe_713_reset = reset;
  assign bc_pe_713_io_ho_input = bc_pe_712_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_713_io_ve_input = bc_pe_681_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_713_io_input_valid = io_input_valid_713; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_713_io_iormac = io_iormac_713; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_714_clock = clock;
  assign bc_pe_714_reset = reset;
  assign bc_pe_714_io_ho_input = bc_pe_713_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_714_io_ve_input = bc_pe_682_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_714_io_input_valid = io_input_valid_714; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_714_io_iormac = io_iormac_714; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_715_clock = clock;
  assign bc_pe_715_reset = reset;
  assign bc_pe_715_io_ho_input = bc_pe_714_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_715_io_ve_input = bc_pe_683_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_715_io_input_valid = io_input_valid_715; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_715_io_iormac = io_iormac_715; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_716_clock = clock;
  assign bc_pe_716_reset = reset;
  assign bc_pe_716_io_ho_input = bc_pe_715_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_716_io_ve_input = bc_pe_684_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_716_io_input_valid = io_input_valid_716; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_716_io_iormac = io_iormac_716; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_717_clock = clock;
  assign bc_pe_717_reset = reset;
  assign bc_pe_717_io_ho_input = bc_pe_716_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_717_io_ve_input = bc_pe_685_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_717_io_input_valid = io_input_valid_717; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_717_io_iormac = io_iormac_717; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_718_clock = clock;
  assign bc_pe_718_reset = reset;
  assign bc_pe_718_io_ho_input = bc_pe_717_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_718_io_ve_input = bc_pe_686_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_718_io_input_valid = io_input_valid_718; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_718_io_iormac = io_iormac_718; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_719_clock = clock;
  assign bc_pe_719_reset = reset;
  assign bc_pe_719_io_ho_input = bc_pe_718_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_719_io_ve_input = bc_pe_687_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_719_io_input_valid = io_input_valid_719; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_719_io_iormac = io_iormac_719; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_720_clock = clock;
  assign bc_pe_720_reset = reset;
  assign bc_pe_720_io_ho_input = bc_pe_719_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_720_io_ve_input = bc_pe_688_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_720_io_input_valid = io_input_valid_720; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_720_io_iormac = io_iormac_720; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_721_clock = clock;
  assign bc_pe_721_reset = reset;
  assign bc_pe_721_io_ho_input = bc_pe_720_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_721_io_ve_input = bc_pe_689_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_721_io_input_valid = io_input_valid_721; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_721_io_iormac = io_iormac_721; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_722_clock = clock;
  assign bc_pe_722_reset = reset;
  assign bc_pe_722_io_ho_input = bc_pe_721_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_722_io_ve_input = bc_pe_690_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_722_io_input_valid = io_input_valid_722; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_722_io_iormac = io_iormac_722; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_723_clock = clock;
  assign bc_pe_723_reset = reset;
  assign bc_pe_723_io_ho_input = bc_pe_722_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_723_io_ve_input = bc_pe_691_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_723_io_input_valid = io_input_valid_723; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_723_io_iormac = io_iormac_723; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_724_clock = clock;
  assign bc_pe_724_reset = reset;
  assign bc_pe_724_io_ho_input = bc_pe_723_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_724_io_ve_input = bc_pe_692_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_724_io_input_valid = io_input_valid_724; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_724_io_iormac = io_iormac_724; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_725_clock = clock;
  assign bc_pe_725_reset = reset;
  assign bc_pe_725_io_ho_input = bc_pe_724_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_725_io_ve_input = bc_pe_693_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_725_io_input_valid = io_input_valid_725; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_725_io_iormac = io_iormac_725; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_726_clock = clock;
  assign bc_pe_726_reset = reset;
  assign bc_pe_726_io_ho_input = bc_pe_725_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_726_io_ve_input = bc_pe_694_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_726_io_input_valid = io_input_valid_726; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_726_io_iormac = io_iormac_726; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_727_clock = clock;
  assign bc_pe_727_reset = reset;
  assign bc_pe_727_io_ho_input = bc_pe_726_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_727_io_ve_input = bc_pe_695_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_727_io_input_valid = io_input_valid_727; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_727_io_iormac = io_iormac_727; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_728_clock = clock;
  assign bc_pe_728_reset = reset;
  assign bc_pe_728_io_ho_input = bc_pe_727_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_728_io_ve_input = bc_pe_696_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_728_io_input_valid = io_input_valid_728; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_728_io_iormac = io_iormac_728; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_729_clock = clock;
  assign bc_pe_729_reset = reset;
  assign bc_pe_729_io_ho_input = bc_pe_728_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_729_io_ve_input = bc_pe_697_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_729_io_input_valid = io_input_valid_729; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_729_io_iormac = io_iormac_729; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_730_clock = clock;
  assign bc_pe_730_reset = reset;
  assign bc_pe_730_io_ho_input = bc_pe_729_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_730_io_ve_input = bc_pe_698_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_730_io_input_valid = io_input_valid_730; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_730_io_iormac = io_iormac_730; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_731_clock = clock;
  assign bc_pe_731_reset = reset;
  assign bc_pe_731_io_ho_input = bc_pe_730_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_731_io_ve_input = bc_pe_699_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_731_io_input_valid = io_input_valid_731; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_731_io_iormac = io_iormac_731; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_732_clock = clock;
  assign bc_pe_732_reset = reset;
  assign bc_pe_732_io_ho_input = bc_pe_731_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_732_io_ve_input = bc_pe_700_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_732_io_input_valid = io_input_valid_732; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_732_io_iormac = io_iormac_732; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_733_clock = clock;
  assign bc_pe_733_reset = reset;
  assign bc_pe_733_io_ho_input = bc_pe_732_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_733_io_ve_input = bc_pe_701_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_733_io_input_valid = io_input_valid_733; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_733_io_iormac = io_iormac_733; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_734_clock = clock;
  assign bc_pe_734_reset = reset;
  assign bc_pe_734_io_ho_input = bc_pe_733_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_734_io_ve_input = bc_pe_702_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_734_io_input_valid = io_input_valid_734; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_734_io_iormac = io_iormac_734; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_735_clock = clock;
  assign bc_pe_735_reset = reset;
  assign bc_pe_735_io_ho_input = bc_pe_734_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_735_io_ve_input = bc_pe_703_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_735_io_input_valid = io_input_valid_735; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_735_io_iormac = io_iormac_735; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_736_clock = clock;
  assign bc_pe_736_reset = reset;
  assign bc_pe_736_io_ho_input = io_x_input_23; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_736_io_ve_input = bc_pe_704_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_736_io_input_valid = io_input_valid_736; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_736_io_iormac = io_iormac_736; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_737_clock = clock;
  assign bc_pe_737_reset = reset;
  assign bc_pe_737_io_ho_input = bc_pe_736_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_737_io_ve_input = bc_pe_705_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_737_io_input_valid = io_input_valid_737; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_737_io_iormac = io_iormac_737; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_738_clock = clock;
  assign bc_pe_738_reset = reset;
  assign bc_pe_738_io_ho_input = bc_pe_737_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_738_io_ve_input = bc_pe_706_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_738_io_input_valid = io_input_valid_738; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_738_io_iormac = io_iormac_738; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_739_clock = clock;
  assign bc_pe_739_reset = reset;
  assign bc_pe_739_io_ho_input = bc_pe_738_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_739_io_ve_input = bc_pe_707_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_739_io_input_valid = io_input_valid_739; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_739_io_iormac = io_iormac_739; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_740_clock = clock;
  assign bc_pe_740_reset = reset;
  assign bc_pe_740_io_ho_input = bc_pe_739_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_740_io_ve_input = bc_pe_708_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_740_io_input_valid = io_input_valid_740; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_740_io_iormac = io_iormac_740; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_741_clock = clock;
  assign bc_pe_741_reset = reset;
  assign bc_pe_741_io_ho_input = bc_pe_740_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_741_io_ve_input = bc_pe_709_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_741_io_input_valid = io_input_valid_741; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_741_io_iormac = io_iormac_741; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_742_clock = clock;
  assign bc_pe_742_reset = reset;
  assign bc_pe_742_io_ho_input = bc_pe_741_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_742_io_ve_input = bc_pe_710_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_742_io_input_valid = io_input_valid_742; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_742_io_iormac = io_iormac_742; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_743_clock = clock;
  assign bc_pe_743_reset = reset;
  assign bc_pe_743_io_ho_input = bc_pe_742_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_743_io_ve_input = bc_pe_711_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_743_io_input_valid = io_input_valid_743; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_743_io_iormac = io_iormac_743; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_744_clock = clock;
  assign bc_pe_744_reset = reset;
  assign bc_pe_744_io_ho_input = bc_pe_743_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_744_io_ve_input = bc_pe_712_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_744_io_input_valid = io_input_valid_744; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_744_io_iormac = io_iormac_744; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_745_clock = clock;
  assign bc_pe_745_reset = reset;
  assign bc_pe_745_io_ho_input = bc_pe_744_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_745_io_ve_input = bc_pe_713_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_745_io_input_valid = io_input_valid_745; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_745_io_iormac = io_iormac_745; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_746_clock = clock;
  assign bc_pe_746_reset = reset;
  assign bc_pe_746_io_ho_input = bc_pe_745_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_746_io_ve_input = bc_pe_714_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_746_io_input_valid = io_input_valid_746; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_746_io_iormac = io_iormac_746; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_747_clock = clock;
  assign bc_pe_747_reset = reset;
  assign bc_pe_747_io_ho_input = bc_pe_746_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_747_io_ve_input = bc_pe_715_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_747_io_input_valid = io_input_valid_747; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_747_io_iormac = io_iormac_747; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_748_clock = clock;
  assign bc_pe_748_reset = reset;
  assign bc_pe_748_io_ho_input = bc_pe_747_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_748_io_ve_input = bc_pe_716_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_748_io_input_valid = io_input_valid_748; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_748_io_iormac = io_iormac_748; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_749_clock = clock;
  assign bc_pe_749_reset = reset;
  assign bc_pe_749_io_ho_input = bc_pe_748_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_749_io_ve_input = bc_pe_717_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_749_io_input_valid = io_input_valid_749; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_749_io_iormac = io_iormac_749; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_750_clock = clock;
  assign bc_pe_750_reset = reset;
  assign bc_pe_750_io_ho_input = bc_pe_749_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_750_io_ve_input = bc_pe_718_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_750_io_input_valid = io_input_valid_750; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_750_io_iormac = io_iormac_750; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_751_clock = clock;
  assign bc_pe_751_reset = reset;
  assign bc_pe_751_io_ho_input = bc_pe_750_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_751_io_ve_input = bc_pe_719_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_751_io_input_valid = io_input_valid_751; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_751_io_iormac = io_iormac_751; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_752_clock = clock;
  assign bc_pe_752_reset = reset;
  assign bc_pe_752_io_ho_input = bc_pe_751_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_752_io_ve_input = bc_pe_720_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_752_io_input_valid = io_input_valid_752; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_752_io_iormac = io_iormac_752; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_753_clock = clock;
  assign bc_pe_753_reset = reset;
  assign bc_pe_753_io_ho_input = bc_pe_752_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_753_io_ve_input = bc_pe_721_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_753_io_input_valid = io_input_valid_753; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_753_io_iormac = io_iormac_753; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_754_clock = clock;
  assign bc_pe_754_reset = reset;
  assign bc_pe_754_io_ho_input = bc_pe_753_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_754_io_ve_input = bc_pe_722_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_754_io_input_valid = io_input_valid_754; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_754_io_iormac = io_iormac_754; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_755_clock = clock;
  assign bc_pe_755_reset = reset;
  assign bc_pe_755_io_ho_input = bc_pe_754_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_755_io_ve_input = bc_pe_723_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_755_io_input_valid = io_input_valid_755; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_755_io_iormac = io_iormac_755; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_756_clock = clock;
  assign bc_pe_756_reset = reset;
  assign bc_pe_756_io_ho_input = bc_pe_755_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_756_io_ve_input = bc_pe_724_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_756_io_input_valid = io_input_valid_756; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_756_io_iormac = io_iormac_756; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_757_clock = clock;
  assign bc_pe_757_reset = reset;
  assign bc_pe_757_io_ho_input = bc_pe_756_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_757_io_ve_input = bc_pe_725_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_757_io_input_valid = io_input_valid_757; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_757_io_iormac = io_iormac_757; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_758_clock = clock;
  assign bc_pe_758_reset = reset;
  assign bc_pe_758_io_ho_input = bc_pe_757_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_758_io_ve_input = bc_pe_726_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_758_io_input_valid = io_input_valid_758; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_758_io_iormac = io_iormac_758; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_759_clock = clock;
  assign bc_pe_759_reset = reset;
  assign bc_pe_759_io_ho_input = bc_pe_758_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_759_io_ve_input = bc_pe_727_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_759_io_input_valid = io_input_valid_759; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_759_io_iormac = io_iormac_759; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_760_clock = clock;
  assign bc_pe_760_reset = reset;
  assign bc_pe_760_io_ho_input = bc_pe_759_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_760_io_ve_input = bc_pe_728_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_760_io_input_valid = io_input_valid_760; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_760_io_iormac = io_iormac_760; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_761_clock = clock;
  assign bc_pe_761_reset = reset;
  assign bc_pe_761_io_ho_input = bc_pe_760_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_761_io_ve_input = bc_pe_729_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_761_io_input_valid = io_input_valid_761; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_761_io_iormac = io_iormac_761; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_762_clock = clock;
  assign bc_pe_762_reset = reset;
  assign bc_pe_762_io_ho_input = bc_pe_761_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_762_io_ve_input = bc_pe_730_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_762_io_input_valid = io_input_valid_762; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_762_io_iormac = io_iormac_762; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_763_clock = clock;
  assign bc_pe_763_reset = reset;
  assign bc_pe_763_io_ho_input = bc_pe_762_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_763_io_ve_input = bc_pe_731_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_763_io_input_valid = io_input_valid_763; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_763_io_iormac = io_iormac_763; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_764_clock = clock;
  assign bc_pe_764_reset = reset;
  assign bc_pe_764_io_ho_input = bc_pe_763_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_764_io_ve_input = bc_pe_732_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_764_io_input_valid = io_input_valid_764; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_764_io_iormac = io_iormac_764; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_765_clock = clock;
  assign bc_pe_765_reset = reset;
  assign bc_pe_765_io_ho_input = bc_pe_764_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_765_io_ve_input = bc_pe_733_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_765_io_input_valid = io_input_valid_765; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_765_io_iormac = io_iormac_765; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_766_clock = clock;
  assign bc_pe_766_reset = reset;
  assign bc_pe_766_io_ho_input = bc_pe_765_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_766_io_ve_input = bc_pe_734_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_766_io_input_valid = io_input_valid_766; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_766_io_iormac = io_iormac_766; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_767_clock = clock;
  assign bc_pe_767_reset = reset;
  assign bc_pe_767_io_ho_input = bc_pe_766_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_767_io_ve_input = bc_pe_735_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_767_io_input_valid = io_input_valid_767; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_767_io_iormac = io_iormac_767; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_768_clock = clock;
  assign bc_pe_768_reset = reset;
  assign bc_pe_768_io_ho_input = io_x_input_24; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_768_io_ve_input = bc_pe_736_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_768_io_input_valid = io_input_valid_768; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_768_io_iormac = io_iormac_768; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_769_clock = clock;
  assign bc_pe_769_reset = reset;
  assign bc_pe_769_io_ho_input = bc_pe_768_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_769_io_ve_input = bc_pe_737_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_769_io_input_valid = io_input_valid_769; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_769_io_iormac = io_iormac_769; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_770_clock = clock;
  assign bc_pe_770_reset = reset;
  assign bc_pe_770_io_ho_input = bc_pe_769_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_770_io_ve_input = bc_pe_738_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_770_io_input_valid = io_input_valid_770; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_770_io_iormac = io_iormac_770; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_771_clock = clock;
  assign bc_pe_771_reset = reset;
  assign bc_pe_771_io_ho_input = bc_pe_770_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_771_io_ve_input = bc_pe_739_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_771_io_input_valid = io_input_valid_771; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_771_io_iormac = io_iormac_771; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_772_clock = clock;
  assign bc_pe_772_reset = reset;
  assign bc_pe_772_io_ho_input = bc_pe_771_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_772_io_ve_input = bc_pe_740_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_772_io_input_valid = io_input_valid_772; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_772_io_iormac = io_iormac_772; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_773_clock = clock;
  assign bc_pe_773_reset = reset;
  assign bc_pe_773_io_ho_input = bc_pe_772_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_773_io_ve_input = bc_pe_741_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_773_io_input_valid = io_input_valid_773; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_773_io_iormac = io_iormac_773; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_774_clock = clock;
  assign bc_pe_774_reset = reset;
  assign bc_pe_774_io_ho_input = bc_pe_773_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_774_io_ve_input = bc_pe_742_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_774_io_input_valid = io_input_valid_774; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_774_io_iormac = io_iormac_774; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_775_clock = clock;
  assign bc_pe_775_reset = reset;
  assign bc_pe_775_io_ho_input = bc_pe_774_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_775_io_ve_input = bc_pe_743_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_775_io_input_valid = io_input_valid_775; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_775_io_iormac = io_iormac_775; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_776_clock = clock;
  assign bc_pe_776_reset = reset;
  assign bc_pe_776_io_ho_input = bc_pe_775_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_776_io_ve_input = bc_pe_744_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_776_io_input_valid = io_input_valid_776; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_776_io_iormac = io_iormac_776; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_777_clock = clock;
  assign bc_pe_777_reset = reset;
  assign bc_pe_777_io_ho_input = bc_pe_776_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_777_io_ve_input = bc_pe_745_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_777_io_input_valid = io_input_valid_777; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_777_io_iormac = io_iormac_777; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_778_clock = clock;
  assign bc_pe_778_reset = reset;
  assign bc_pe_778_io_ho_input = bc_pe_777_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_778_io_ve_input = bc_pe_746_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_778_io_input_valid = io_input_valid_778; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_778_io_iormac = io_iormac_778; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_779_clock = clock;
  assign bc_pe_779_reset = reset;
  assign bc_pe_779_io_ho_input = bc_pe_778_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_779_io_ve_input = bc_pe_747_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_779_io_input_valid = io_input_valid_779; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_779_io_iormac = io_iormac_779; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_780_clock = clock;
  assign bc_pe_780_reset = reset;
  assign bc_pe_780_io_ho_input = bc_pe_779_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_780_io_ve_input = bc_pe_748_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_780_io_input_valid = io_input_valid_780; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_780_io_iormac = io_iormac_780; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_781_clock = clock;
  assign bc_pe_781_reset = reset;
  assign bc_pe_781_io_ho_input = bc_pe_780_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_781_io_ve_input = bc_pe_749_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_781_io_input_valid = io_input_valid_781; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_781_io_iormac = io_iormac_781; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_782_clock = clock;
  assign bc_pe_782_reset = reset;
  assign bc_pe_782_io_ho_input = bc_pe_781_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_782_io_ve_input = bc_pe_750_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_782_io_input_valid = io_input_valid_782; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_782_io_iormac = io_iormac_782; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_783_clock = clock;
  assign bc_pe_783_reset = reset;
  assign bc_pe_783_io_ho_input = bc_pe_782_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_783_io_ve_input = bc_pe_751_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_783_io_input_valid = io_input_valid_783; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_783_io_iormac = io_iormac_783; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_784_clock = clock;
  assign bc_pe_784_reset = reset;
  assign bc_pe_784_io_ho_input = bc_pe_783_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_784_io_ve_input = bc_pe_752_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_784_io_input_valid = io_input_valid_784; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_784_io_iormac = io_iormac_784; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_785_clock = clock;
  assign bc_pe_785_reset = reset;
  assign bc_pe_785_io_ho_input = bc_pe_784_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_785_io_ve_input = bc_pe_753_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_785_io_input_valid = io_input_valid_785; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_785_io_iormac = io_iormac_785; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_786_clock = clock;
  assign bc_pe_786_reset = reset;
  assign bc_pe_786_io_ho_input = bc_pe_785_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_786_io_ve_input = bc_pe_754_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_786_io_input_valid = io_input_valid_786; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_786_io_iormac = io_iormac_786; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_787_clock = clock;
  assign bc_pe_787_reset = reset;
  assign bc_pe_787_io_ho_input = bc_pe_786_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_787_io_ve_input = bc_pe_755_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_787_io_input_valid = io_input_valid_787; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_787_io_iormac = io_iormac_787; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_788_clock = clock;
  assign bc_pe_788_reset = reset;
  assign bc_pe_788_io_ho_input = bc_pe_787_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_788_io_ve_input = bc_pe_756_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_788_io_input_valid = io_input_valid_788; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_788_io_iormac = io_iormac_788; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_789_clock = clock;
  assign bc_pe_789_reset = reset;
  assign bc_pe_789_io_ho_input = bc_pe_788_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_789_io_ve_input = bc_pe_757_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_789_io_input_valid = io_input_valid_789; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_789_io_iormac = io_iormac_789; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_790_clock = clock;
  assign bc_pe_790_reset = reset;
  assign bc_pe_790_io_ho_input = bc_pe_789_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_790_io_ve_input = bc_pe_758_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_790_io_input_valid = io_input_valid_790; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_790_io_iormac = io_iormac_790; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_791_clock = clock;
  assign bc_pe_791_reset = reset;
  assign bc_pe_791_io_ho_input = bc_pe_790_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_791_io_ve_input = bc_pe_759_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_791_io_input_valid = io_input_valid_791; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_791_io_iormac = io_iormac_791; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_792_clock = clock;
  assign bc_pe_792_reset = reset;
  assign bc_pe_792_io_ho_input = bc_pe_791_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_792_io_ve_input = bc_pe_760_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_792_io_input_valid = io_input_valid_792; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_792_io_iormac = io_iormac_792; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_793_clock = clock;
  assign bc_pe_793_reset = reset;
  assign bc_pe_793_io_ho_input = bc_pe_792_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_793_io_ve_input = bc_pe_761_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_793_io_input_valid = io_input_valid_793; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_793_io_iormac = io_iormac_793; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_794_clock = clock;
  assign bc_pe_794_reset = reset;
  assign bc_pe_794_io_ho_input = bc_pe_793_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_794_io_ve_input = bc_pe_762_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_794_io_input_valid = io_input_valid_794; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_794_io_iormac = io_iormac_794; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_795_clock = clock;
  assign bc_pe_795_reset = reset;
  assign bc_pe_795_io_ho_input = bc_pe_794_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_795_io_ve_input = bc_pe_763_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_795_io_input_valid = io_input_valid_795; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_795_io_iormac = io_iormac_795; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_796_clock = clock;
  assign bc_pe_796_reset = reset;
  assign bc_pe_796_io_ho_input = bc_pe_795_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_796_io_ve_input = bc_pe_764_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_796_io_input_valid = io_input_valid_796; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_796_io_iormac = io_iormac_796; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_797_clock = clock;
  assign bc_pe_797_reset = reset;
  assign bc_pe_797_io_ho_input = bc_pe_796_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_797_io_ve_input = bc_pe_765_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_797_io_input_valid = io_input_valid_797; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_797_io_iormac = io_iormac_797; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_798_clock = clock;
  assign bc_pe_798_reset = reset;
  assign bc_pe_798_io_ho_input = bc_pe_797_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_798_io_ve_input = bc_pe_766_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_798_io_input_valid = io_input_valid_798; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_798_io_iormac = io_iormac_798; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_799_clock = clock;
  assign bc_pe_799_reset = reset;
  assign bc_pe_799_io_ho_input = bc_pe_798_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_799_io_ve_input = bc_pe_767_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_799_io_input_valid = io_input_valid_799; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_799_io_iormac = io_iormac_799; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_800_clock = clock;
  assign bc_pe_800_reset = reset;
  assign bc_pe_800_io_ho_input = io_x_input_25; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_800_io_ve_input = bc_pe_768_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_800_io_input_valid = io_input_valid_800; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_800_io_iormac = io_iormac_800; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_801_clock = clock;
  assign bc_pe_801_reset = reset;
  assign bc_pe_801_io_ho_input = bc_pe_800_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_801_io_ve_input = bc_pe_769_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_801_io_input_valid = io_input_valid_801; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_801_io_iormac = io_iormac_801; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_802_clock = clock;
  assign bc_pe_802_reset = reset;
  assign bc_pe_802_io_ho_input = bc_pe_801_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_802_io_ve_input = bc_pe_770_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_802_io_input_valid = io_input_valid_802; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_802_io_iormac = io_iormac_802; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_803_clock = clock;
  assign bc_pe_803_reset = reset;
  assign bc_pe_803_io_ho_input = bc_pe_802_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_803_io_ve_input = bc_pe_771_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_803_io_input_valid = io_input_valid_803; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_803_io_iormac = io_iormac_803; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_804_clock = clock;
  assign bc_pe_804_reset = reset;
  assign bc_pe_804_io_ho_input = bc_pe_803_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_804_io_ve_input = bc_pe_772_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_804_io_input_valid = io_input_valid_804; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_804_io_iormac = io_iormac_804; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_805_clock = clock;
  assign bc_pe_805_reset = reset;
  assign bc_pe_805_io_ho_input = bc_pe_804_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_805_io_ve_input = bc_pe_773_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_805_io_input_valid = io_input_valid_805; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_805_io_iormac = io_iormac_805; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_806_clock = clock;
  assign bc_pe_806_reset = reset;
  assign bc_pe_806_io_ho_input = bc_pe_805_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_806_io_ve_input = bc_pe_774_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_806_io_input_valid = io_input_valid_806; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_806_io_iormac = io_iormac_806; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_807_clock = clock;
  assign bc_pe_807_reset = reset;
  assign bc_pe_807_io_ho_input = bc_pe_806_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_807_io_ve_input = bc_pe_775_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_807_io_input_valid = io_input_valid_807; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_807_io_iormac = io_iormac_807; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_808_clock = clock;
  assign bc_pe_808_reset = reset;
  assign bc_pe_808_io_ho_input = bc_pe_807_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_808_io_ve_input = bc_pe_776_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_808_io_input_valid = io_input_valid_808; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_808_io_iormac = io_iormac_808; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_809_clock = clock;
  assign bc_pe_809_reset = reset;
  assign bc_pe_809_io_ho_input = bc_pe_808_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_809_io_ve_input = bc_pe_777_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_809_io_input_valid = io_input_valid_809; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_809_io_iormac = io_iormac_809; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_810_clock = clock;
  assign bc_pe_810_reset = reset;
  assign bc_pe_810_io_ho_input = bc_pe_809_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_810_io_ve_input = bc_pe_778_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_810_io_input_valid = io_input_valid_810; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_810_io_iormac = io_iormac_810; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_811_clock = clock;
  assign bc_pe_811_reset = reset;
  assign bc_pe_811_io_ho_input = bc_pe_810_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_811_io_ve_input = bc_pe_779_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_811_io_input_valid = io_input_valid_811; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_811_io_iormac = io_iormac_811; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_812_clock = clock;
  assign bc_pe_812_reset = reset;
  assign bc_pe_812_io_ho_input = bc_pe_811_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_812_io_ve_input = bc_pe_780_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_812_io_input_valid = io_input_valid_812; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_812_io_iormac = io_iormac_812; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_813_clock = clock;
  assign bc_pe_813_reset = reset;
  assign bc_pe_813_io_ho_input = bc_pe_812_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_813_io_ve_input = bc_pe_781_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_813_io_input_valid = io_input_valid_813; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_813_io_iormac = io_iormac_813; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_814_clock = clock;
  assign bc_pe_814_reset = reset;
  assign bc_pe_814_io_ho_input = bc_pe_813_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_814_io_ve_input = bc_pe_782_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_814_io_input_valid = io_input_valid_814; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_814_io_iormac = io_iormac_814; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_815_clock = clock;
  assign bc_pe_815_reset = reset;
  assign bc_pe_815_io_ho_input = bc_pe_814_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_815_io_ve_input = bc_pe_783_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_815_io_input_valid = io_input_valid_815; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_815_io_iormac = io_iormac_815; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_816_clock = clock;
  assign bc_pe_816_reset = reset;
  assign bc_pe_816_io_ho_input = bc_pe_815_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_816_io_ve_input = bc_pe_784_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_816_io_input_valid = io_input_valid_816; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_816_io_iormac = io_iormac_816; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_817_clock = clock;
  assign bc_pe_817_reset = reset;
  assign bc_pe_817_io_ho_input = bc_pe_816_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_817_io_ve_input = bc_pe_785_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_817_io_input_valid = io_input_valid_817; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_817_io_iormac = io_iormac_817; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_818_clock = clock;
  assign bc_pe_818_reset = reset;
  assign bc_pe_818_io_ho_input = bc_pe_817_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_818_io_ve_input = bc_pe_786_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_818_io_input_valid = io_input_valid_818; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_818_io_iormac = io_iormac_818; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_819_clock = clock;
  assign bc_pe_819_reset = reset;
  assign bc_pe_819_io_ho_input = bc_pe_818_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_819_io_ve_input = bc_pe_787_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_819_io_input_valid = io_input_valid_819; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_819_io_iormac = io_iormac_819; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_820_clock = clock;
  assign bc_pe_820_reset = reset;
  assign bc_pe_820_io_ho_input = bc_pe_819_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_820_io_ve_input = bc_pe_788_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_820_io_input_valid = io_input_valid_820; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_820_io_iormac = io_iormac_820; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_821_clock = clock;
  assign bc_pe_821_reset = reset;
  assign bc_pe_821_io_ho_input = bc_pe_820_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_821_io_ve_input = bc_pe_789_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_821_io_input_valid = io_input_valid_821; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_821_io_iormac = io_iormac_821; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_822_clock = clock;
  assign bc_pe_822_reset = reset;
  assign bc_pe_822_io_ho_input = bc_pe_821_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_822_io_ve_input = bc_pe_790_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_822_io_input_valid = io_input_valid_822; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_822_io_iormac = io_iormac_822; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_823_clock = clock;
  assign bc_pe_823_reset = reset;
  assign bc_pe_823_io_ho_input = bc_pe_822_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_823_io_ve_input = bc_pe_791_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_823_io_input_valid = io_input_valid_823; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_823_io_iormac = io_iormac_823; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_824_clock = clock;
  assign bc_pe_824_reset = reset;
  assign bc_pe_824_io_ho_input = bc_pe_823_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_824_io_ve_input = bc_pe_792_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_824_io_input_valid = io_input_valid_824; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_824_io_iormac = io_iormac_824; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_825_clock = clock;
  assign bc_pe_825_reset = reset;
  assign bc_pe_825_io_ho_input = bc_pe_824_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_825_io_ve_input = bc_pe_793_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_825_io_input_valid = io_input_valid_825; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_825_io_iormac = io_iormac_825; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_826_clock = clock;
  assign bc_pe_826_reset = reset;
  assign bc_pe_826_io_ho_input = bc_pe_825_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_826_io_ve_input = bc_pe_794_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_826_io_input_valid = io_input_valid_826; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_826_io_iormac = io_iormac_826; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_827_clock = clock;
  assign bc_pe_827_reset = reset;
  assign bc_pe_827_io_ho_input = bc_pe_826_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_827_io_ve_input = bc_pe_795_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_827_io_input_valid = io_input_valid_827; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_827_io_iormac = io_iormac_827; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_828_clock = clock;
  assign bc_pe_828_reset = reset;
  assign bc_pe_828_io_ho_input = bc_pe_827_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_828_io_ve_input = bc_pe_796_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_828_io_input_valid = io_input_valid_828; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_828_io_iormac = io_iormac_828; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_829_clock = clock;
  assign bc_pe_829_reset = reset;
  assign bc_pe_829_io_ho_input = bc_pe_828_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_829_io_ve_input = bc_pe_797_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_829_io_input_valid = io_input_valid_829; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_829_io_iormac = io_iormac_829; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_830_clock = clock;
  assign bc_pe_830_reset = reset;
  assign bc_pe_830_io_ho_input = bc_pe_829_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_830_io_ve_input = bc_pe_798_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_830_io_input_valid = io_input_valid_830; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_830_io_iormac = io_iormac_830; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_831_clock = clock;
  assign bc_pe_831_reset = reset;
  assign bc_pe_831_io_ho_input = bc_pe_830_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_831_io_ve_input = bc_pe_799_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_831_io_input_valid = io_input_valid_831; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_831_io_iormac = io_iormac_831; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_832_clock = clock;
  assign bc_pe_832_reset = reset;
  assign bc_pe_832_io_ho_input = io_x_input_26; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_832_io_ve_input = bc_pe_800_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_832_io_input_valid = io_input_valid_832; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_832_io_iormac = io_iormac_832; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_833_clock = clock;
  assign bc_pe_833_reset = reset;
  assign bc_pe_833_io_ho_input = bc_pe_832_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_833_io_ve_input = bc_pe_801_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_833_io_input_valid = io_input_valid_833; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_833_io_iormac = io_iormac_833; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_834_clock = clock;
  assign bc_pe_834_reset = reset;
  assign bc_pe_834_io_ho_input = bc_pe_833_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_834_io_ve_input = bc_pe_802_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_834_io_input_valid = io_input_valid_834; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_834_io_iormac = io_iormac_834; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_835_clock = clock;
  assign bc_pe_835_reset = reset;
  assign bc_pe_835_io_ho_input = bc_pe_834_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_835_io_ve_input = bc_pe_803_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_835_io_input_valid = io_input_valid_835; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_835_io_iormac = io_iormac_835; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_836_clock = clock;
  assign bc_pe_836_reset = reset;
  assign bc_pe_836_io_ho_input = bc_pe_835_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_836_io_ve_input = bc_pe_804_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_836_io_input_valid = io_input_valid_836; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_836_io_iormac = io_iormac_836; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_837_clock = clock;
  assign bc_pe_837_reset = reset;
  assign bc_pe_837_io_ho_input = bc_pe_836_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_837_io_ve_input = bc_pe_805_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_837_io_input_valid = io_input_valid_837; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_837_io_iormac = io_iormac_837; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_838_clock = clock;
  assign bc_pe_838_reset = reset;
  assign bc_pe_838_io_ho_input = bc_pe_837_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_838_io_ve_input = bc_pe_806_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_838_io_input_valid = io_input_valid_838; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_838_io_iormac = io_iormac_838; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_839_clock = clock;
  assign bc_pe_839_reset = reset;
  assign bc_pe_839_io_ho_input = bc_pe_838_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_839_io_ve_input = bc_pe_807_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_839_io_input_valid = io_input_valid_839; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_839_io_iormac = io_iormac_839; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_840_clock = clock;
  assign bc_pe_840_reset = reset;
  assign bc_pe_840_io_ho_input = bc_pe_839_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_840_io_ve_input = bc_pe_808_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_840_io_input_valid = io_input_valid_840; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_840_io_iormac = io_iormac_840; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_841_clock = clock;
  assign bc_pe_841_reset = reset;
  assign bc_pe_841_io_ho_input = bc_pe_840_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_841_io_ve_input = bc_pe_809_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_841_io_input_valid = io_input_valid_841; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_841_io_iormac = io_iormac_841; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_842_clock = clock;
  assign bc_pe_842_reset = reset;
  assign bc_pe_842_io_ho_input = bc_pe_841_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_842_io_ve_input = bc_pe_810_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_842_io_input_valid = io_input_valid_842; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_842_io_iormac = io_iormac_842; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_843_clock = clock;
  assign bc_pe_843_reset = reset;
  assign bc_pe_843_io_ho_input = bc_pe_842_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_843_io_ve_input = bc_pe_811_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_843_io_input_valid = io_input_valid_843; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_843_io_iormac = io_iormac_843; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_844_clock = clock;
  assign bc_pe_844_reset = reset;
  assign bc_pe_844_io_ho_input = bc_pe_843_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_844_io_ve_input = bc_pe_812_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_844_io_input_valid = io_input_valid_844; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_844_io_iormac = io_iormac_844; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_845_clock = clock;
  assign bc_pe_845_reset = reset;
  assign bc_pe_845_io_ho_input = bc_pe_844_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_845_io_ve_input = bc_pe_813_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_845_io_input_valid = io_input_valid_845; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_845_io_iormac = io_iormac_845; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_846_clock = clock;
  assign bc_pe_846_reset = reset;
  assign bc_pe_846_io_ho_input = bc_pe_845_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_846_io_ve_input = bc_pe_814_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_846_io_input_valid = io_input_valid_846; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_846_io_iormac = io_iormac_846; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_847_clock = clock;
  assign bc_pe_847_reset = reset;
  assign bc_pe_847_io_ho_input = bc_pe_846_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_847_io_ve_input = bc_pe_815_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_847_io_input_valid = io_input_valid_847; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_847_io_iormac = io_iormac_847; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_848_clock = clock;
  assign bc_pe_848_reset = reset;
  assign bc_pe_848_io_ho_input = bc_pe_847_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_848_io_ve_input = bc_pe_816_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_848_io_input_valid = io_input_valid_848; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_848_io_iormac = io_iormac_848; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_849_clock = clock;
  assign bc_pe_849_reset = reset;
  assign bc_pe_849_io_ho_input = bc_pe_848_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_849_io_ve_input = bc_pe_817_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_849_io_input_valid = io_input_valid_849; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_849_io_iormac = io_iormac_849; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_850_clock = clock;
  assign bc_pe_850_reset = reset;
  assign bc_pe_850_io_ho_input = bc_pe_849_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_850_io_ve_input = bc_pe_818_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_850_io_input_valid = io_input_valid_850; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_850_io_iormac = io_iormac_850; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_851_clock = clock;
  assign bc_pe_851_reset = reset;
  assign bc_pe_851_io_ho_input = bc_pe_850_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_851_io_ve_input = bc_pe_819_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_851_io_input_valid = io_input_valid_851; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_851_io_iormac = io_iormac_851; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_852_clock = clock;
  assign bc_pe_852_reset = reset;
  assign bc_pe_852_io_ho_input = bc_pe_851_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_852_io_ve_input = bc_pe_820_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_852_io_input_valid = io_input_valid_852; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_852_io_iormac = io_iormac_852; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_853_clock = clock;
  assign bc_pe_853_reset = reset;
  assign bc_pe_853_io_ho_input = bc_pe_852_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_853_io_ve_input = bc_pe_821_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_853_io_input_valid = io_input_valid_853; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_853_io_iormac = io_iormac_853; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_854_clock = clock;
  assign bc_pe_854_reset = reset;
  assign bc_pe_854_io_ho_input = bc_pe_853_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_854_io_ve_input = bc_pe_822_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_854_io_input_valid = io_input_valid_854; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_854_io_iormac = io_iormac_854; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_855_clock = clock;
  assign bc_pe_855_reset = reset;
  assign bc_pe_855_io_ho_input = bc_pe_854_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_855_io_ve_input = bc_pe_823_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_855_io_input_valid = io_input_valid_855; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_855_io_iormac = io_iormac_855; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_856_clock = clock;
  assign bc_pe_856_reset = reset;
  assign bc_pe_856_io_ho_input = bc_pe_855_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_856_io_ve_input = bc_pe_824_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_856_io_input_valid = io_input_valid_856; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_856_io_iormac = io_iormac_856; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_857_clock = clock;
  assign bc_pe_857_reset = reset;
  assign bc_pe_857_io_ho_input = bc_pe_856_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_857_io_ve_input = bc_pe_825_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_857_io_input_valid = io_input_valid_857; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_857_io_iormac = io_iormac_857; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_858_clock = clock;
  assign bc_pe_858_reset = reset;
  assign bc_pe_858_io_ho_input = bc_pe_857_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_858_io_ve_input = bc_pe_826_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_858_io_input_valid = io_input_valid_858; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_858_io_iormac = io_iormac_858; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_859_clock = clock;
  assign bc_pe_859_reset = reset;
  assign bc_pe_859_io_ho_input = bc_pe_858_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_859_io_ve_input = bc_pe_827_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_859_io_input_valid = io_input_valid_859; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_859_io_iormac = io_iormac_859; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_860_clock = clock;
  assign bc_pe_860_reset = reset;
  assign bc_pe_860_io_ho_input = bc_pe_859_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_860_io_ve_input = bc_pe_828_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_860_io_input_valid = io_input_valid_860; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_860_io_iormac = io_iormac_860; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_861_clock = clock;
  assign bc_pe_861_reset = reset;
  assign bc_pe_861_io_ho_input = bc_pe_860_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_861_io_ve_input = bc_pe_829_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_861_io_input_valid = io_input_valid_861; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_861_io_iormac = io_iormac_861; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_862_clock = clock;
  assign bc_pe_862_reset = reset;
  assign bc_pe_862_io_ho_input = bc_pe_861_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_862_io_ve_input = bc_pe_830_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_862_io_input_valid = io_input_valid_862; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_862_io_iormac = io_iormac_862; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_863_clock = clock;
  assign bc_pe_863_reset = reset;
  assign bc_pe_863_io_ho_input = bc_pe_862_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_863_io_ve_input = bc_pe_831_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_863_io_input_valid = io_input_valid_863; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_863_io_iormac = io_iormac_863; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_864_clock = clock;
  assign bc_pe_864_reset = reset;
  assign bc_pe_864_io_ho_input = io_x_input_27; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_864_io_ve_input = bc_pe_832_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_864_io_input_valid = io_input_valid_864; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_864_io_iormac = io_iormac_864; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_865_clock = clock;
  assign bc_pe_865_reset = reset;
  assign bc_pe_865_io_ho_input = bc_pe_864_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_865_io_ve_input = bc_pe_833_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_865_io_input_valid = io_input_valid_865; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_865_io_iormac = io_iormac_865; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_866_clock = clock;
  assign bc_pe_866_reset = reset;
  assign bc_pe_866_io_ho_input = bc_pe_865_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_866_io_ve_input = bc_pe_834_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_866_io_input_valid = io_input_valid_866; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_866_io_iormac = io_iormac_866; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_867_clock = clock;
  assign bc_pe_867_reset = reset;
  assign bc_pe_867_io_ho_input = bc_pe_866_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_867_io_ve_input = bc_pe_835_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_867_io_input_valid = io_input_valid_867; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_867_io_iormac = io_iormac_867; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_868_clock = clock;
  assign bc_pe_868_reset = reset;
  assign bc_pe_868_io_ho_input = bc_pe_867_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_868_io_ve_input = bc_pe_836_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_868_io_input_valid = io_input_valid_868; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_868_io_iormac = io_iormac_868; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_869_clock = clock;
  assign bc_pe_869_reset = reset;
  assign bc_pe_869_io_ho_input = bc_pe_868_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_869_io_ve_input = bc_pe_837_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_869_io_input_valid = io_input_valid_869; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_869_io_iormac = io_iormac_869; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_870_clock = clock;
  assign bc_pe_870_reset = reset;
  assign bc_pe_870_io_ho_input = bc_pe_869_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_870_io_ve_input = bc_pe_838_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_870_io_input_valid = io_input_valid_870; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_870_io_iormac = io_iormac_870; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_871_clock = clock;
  assign bc_pe_871_reset = reset;
  assign bc_pe_871_io_ho_input = bc_pe_870_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_871_io_ve_input = bc_pe_839_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_871_io_input_valid = io_input_valid_871; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_871_io_iormac = io_iormac_871; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_872_clock = clock;
  assign bc_pe_872_reset = reset;
  assign bc_pe_872_io_ho_input = bc_pe_871_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_872_io_ve_input = bc_pe_840_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_872_io_input_valid = io_input_valid_872; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_872_io_iormac = io_iormac_872; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_873_clock = clock;
  assign bc_pe_873_reset = reset;
  assign bc_pe_873_io_ho_input = bc_pe_872_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_873_io_ve_input = bc_pe_841_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_873_io_input_valid = io_input_valid_873; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_873_io_iormac = io_iormac_873; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_874_clock = clock;
  assign bc_pe_874_reset = reset;
  assign bc_pe_874_io_ho_input = bc_pe_873_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_874_io_ve_input = bc_pe_842_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_874_io_input_valid = io_input_valid_874; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_874_io_iormac = io_iormac_874; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_875_clock = clock;
  assign bc_pe_875_reset = reset;
  assign bc_pe_875_io_ho_input = bc_pe_874_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_875_io_ve_input = bc_pe_843_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_875_io_input_valid = io_input_valid_875; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_875_io_iormac = io_iormac_875; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_876_clock = clock;
  assign bc_pe_876_reset = reset;
  assign bc_pe_876_io_ho_input = bc_pe_875_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_876_io_ve_input = bc_pe_844_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_876_io_input_valid = io_input_valid_876; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_876_io_iormac = io_iormac_876; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_877_clock = clock;
  assign bc_pe_877_reset = reset;
  assign bc_pe_877_io_ho_input = bc_pe_876_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_877_io_ve_input = bc_pe_845_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_877_io_input_valid = io_input_valid_877; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_877_io_iormac = io_iormac_877; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_878_clock = clock;
  assign bc_pe_878_reset = reset;
  assign bc_pe_878_io_ho_input = bc_pe_877_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_878_io_ve_input = bc_pe_846_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_878_io_input_valid = io_input_valid_878; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_878_io_iormac = io_iormac_878; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_879_clock = clock;
  assign bc_pe_879_reset = reset;
  assign bc_pe_879_io_ho_input = bc_pe_878_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_879_io_ve_input = bc_pe_847_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_879_io_input_valid = io_input_valid_879; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_879_io_iormac = io_iormac_879; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_880_clock = clock;
  assign bc_pe_880_reset = reset;
  assign bc_pe_880_io_ho_input = bc_pe_879_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_880_io_ve_input = bc_pe_848_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_880_io_input_valid = io_input_valid_880; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_880_io_iormac = io_iormac_880; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_881_clock = clock;
  assign bc_pe_881_reset = reset;
  assign bc_pe_881_io_ho_input = bc_pe_880_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_881_io_ve_input = bc_pe_849_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_881_io_input_valid = io_input_valid_881; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_881_io_iormac = io_iormac_881; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_882_clock = clock;
  assign bc_pe_882_reset = reset;
  assign bc_pe_882_io_ho_input = bc_pe_881_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_882_io_ve_input = bc_pe_850_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_882_io_input_valid = io_input_valid_882; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_882_io_iormac = io_iormac_882; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_883_clock = clock;
  assign bc_pe_883_reset = reset;
  assign bc_pe_883_io_ho_input = bc_pe_882_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_883_io_ve_input = bc_pe_851_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_883_io_input_valid = io_input_valid_883; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_883_io_iormac = io_iormac_883; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_884_clock = clock;
  assign bc_pe_884_reset = reset;
  assign bc_pe_884_io_ho_input = bc_pe_883_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_884_io_ve_input = bc_pe_852_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_884_io_input_valid = io_input_valid_884; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_884_io_iormac = io_iormac_884; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_885_clock = clock;
  assign bc_pe_885_reset = reset;
  assign bc_pe_885_io_ho_input = bc_pe_884_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_885_io_ve_input = bc_pe_853_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_885_io_input_valid = io_input_valid_885; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_885_io_iormac = io_iormac_885; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_886_clock = clock;
  assign bc_pe_886_reset = reset;
  assign bc_pe_886_io_ho_input = bc_pe_885_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_886_io_ve_input = bc_pe_854_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_886_io_input_valid = io_input_valid_886; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_886_io_iormac = io_iormac_886; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_887_clock = clock;
  assign bc_pe_887_reset = reset;
  assign bc_pe_887_io_ho_input = bc_pe_886_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_887_io_ve_input = bc_pe_855_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_887_io_input_valid = io_input_valid_887; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_887_io_iormac = io_iormac_887; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_888_clock = clock;
  assign bc_pe_888_reset = reset;
  assign bc_pe_888_io_ho_input = bc_pe_887_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_888_io_ve_input = bc_pe_856_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_888_io_input_valid = io_input_valid_888; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_888_io_iormac = io_iormac_888; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_889_clock = clock;
  assign bc_pe_889_reset = reset;
  assign bc_pe_889_io_ho_input = bc_pe_888_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_889_io_ve_input = bc_pe_857_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_889_io_input_valid = io_input_valid_889; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_889_io_iormac = io_iormac_889; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_890_clock = clock;
  assign bc_pe_890_reset = reset;
  assign bc_pe_890_io_ho_input = bc_pe_889_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_890_io_ve_input = bc_pe_858_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_890_io_input_valid = io_input_valid_890; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_890_io_iormac = io_iormac_890; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_891_clock = clock;
  assign bc_pe_891_reset = reset;
  assign bc_pe_891_io_ho_input = bc_pe_890_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_891_io_ve_input = bc_pe_859_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_891_io_input_valid = io_input_valid_891; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_891_io_iormac = io_iormac_891; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_892_clock = clock;
  assign bc_pe_892_reset = reset;
  assign bc_pe_892_io_ho_input = bc_pe_891_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_892_io_ve_input = bc_pe_860_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_892_io_input_valid = io_input_valid_892; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_892_io_iormac = io_iormac_892; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_893_clock = clock;
  assign bc_pe_893_reset = reset;
  assign bc_pe_893_io_ho_input = bc_pe_892_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_893_io_ve_input = bc_pe_861_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_893_io_input_valid = io_input_valid_893; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_893_io_iormac = io_iormac_893; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_894_clock = clock;
  assign bc_pe_894_reset = reset;
  assign bc_pe_894_io_ho_input = bc_pe_893_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_894_io_ve_input = bc_pe_862_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_894_io_input_valid = io_input_valid_894; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_894_io_iormac = io_iormac_894; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_895_clock = clock;
  assign bc_pe_895_reset = reset;
  assign bc_pe_895_io_ho_input = bc_pe_894_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_895_io_ve_input = bc_pe_863_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_895_io_input_valid = io_input_valid_895; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_895_io_iormac = io_iormac_895; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_896_clock = clock;
  assign bc_pe_896_reset = reset;
  assign bc_pe_896_io_ho_input = io_x_input_28; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_896_io_ve_input = bc_pe_864_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_896_io_input_valid = io_input_valid_896; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_896_io_iormac = io_iormac_896; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_897_clock = clock;
  assign bc_pe_897_reset = reset;
  assign bc_pe_897_io_ho_input = bc_pe_896_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_897_io_ve_input = bc_pe_865_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_897_io_input_valid = io_input_valid_897; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_897_io_iormac = io_iormac_897; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_898_clock = clock;
  assign bc_pe_898_reset = reset;
  assign bc_pe_898_io_ho_input = bc_pe_897_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_898_io_ve_input = bc_pe_866_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_898_io_input_valid = io_input_valid_898; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_898_io_iormac = io_iormac_898; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_899_clock = clock;
  assign bc_pe_899_reset = reset;
  assign bc_pe_899_io_ho_input = bc_pe_898_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_899_io_ve_input = bc_pe_867_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_899_io_input_valid = io_input_valid_899; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_899_io_iormac = io_iormac_899; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_900_clock = clock;
  assign bc_pe_900_reset = reset;
  assign bc_pe_900_io_ho_input = bc_pe_899_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_900_io_ve_input = bc_pe_868_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_900_io_input_valid = io_input_valid_900; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_900_io_iormac = io_iormac_900; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_901_clock = clock;
  assign bc_pe_901_reset = reset;
  assign bc_pe_901_io_ho_input = bc_pe_900_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_901_io_ve_input = bc_pe_869_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_901_io_input_valid = io_input_valid_901; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_901_io_iormac = io_iormac_901; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_902_clock = clock;
  assign bc_pe_902_reset = reset;
  assign bc_pe_902_io_ho_input = bc_pe_901_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_902_io_ve_input = bc_pe_870_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_902_io_input_valid = io_input_valid_902; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_902_io_iormac = io_iormac_902; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_903_clock = clock;
  assign bc_pe_903_reset = reset;
  assign bc_pe_903_io_ho_input = bc_pe_902_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_903_io_ve_input = bc_pe_871_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_903_io_input_valid = io_input_valid_903; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_903_io_iormac = io_iormac_903; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_904_clock = clock;
  assign bc_pe_904_reset = reset;
  assign bc_pe_904_io_ho_input = bc_pe_903_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_904_io_ve_input = bc_pe_872_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_904_io_input_valid = io_input_valid_904; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_904_io_iormac = io_iormac_904; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_905_clock = clock;
  assign bc_pe_905_reset = reset;
  assign bc_pe_905_io_ho_input = bc_pe_904_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_905_io_ve_input = bc_pe_873_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_905_io_input_valid = io_input_valid_905; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_905_io_iormac = io_iormac_905; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_906_clock = clock;
  assign bc_pe_906_reset = reset;
  assign bc_pe_906_io_ho_input = bc_pe_905_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_906_io_ve_input = bc_pe_874_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_906_io_input_valid = io_input_valid_906; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_906_io_iormac = io_iormac_906; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_907_clock = clock;
  assign bc_pe_907_reset = reset;
  assign bc_pe_907_io_ho_input = bc_pe_906_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_907_io_ve_input = bc_pe_875_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_907_io_input_valid = io_input_valid_907; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_907_io_iormac = io_iormac_907; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_908_clock = clock;
  assign bc_pe_908_reset = reset;
  assign bc_pe_908_io_ho_input = bc_pe_907_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_908_io_ve_input = bc_pe_876_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_908_io_input_valid = io_input_valid_908; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_908_io_iormac = io_iormac_908; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_909_clock = clock;
  assign bc_pe_909_reset = reset;
  assign bc_pe_909_io_ho_input = bc_pe_908_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_909_io_ve_input = bc_pe_877_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_909_io_input_valid = io_input_valid_909; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_909_io_iormac = io_iormac_909; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_910_clock = clock;
  assign bc_pe_910_reset = reset;
  assign bc_pe_910_io_ho_input = bc_pe_909_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_910_io_ve_input = bc_pe_878_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_910_io_input_valid = io_input_valid_910; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_910_io_iormac = io_iormac_910; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_911_clock = clock;
  assign bc_pe_911_reset = reset;
  assign bc_pe_911_io_ho_input = bc_pe_910_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_911_io_ve_input = bc_pe_879_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_911_io_input_valid = io_input_valid_911; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_911_io_iormac = io_iormac_911; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_912_clock = clock;
  assign bc_pe_912_reset = reset;
  assign bc_pe_912_io_ho_input = bc_pe_911_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_912_io_ve_input = bc_pe_880_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_912_io_input_valid = io_input_valid_912; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_912_io_iormac = io_iormac_912; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_913_clock = clock;
  assign bc_pe_913_reset = reset;
  assign bc_pe_913_io_ho_input = bc_pe_912_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_913_io_ve_input = bc_pe_881_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_913_io_input_valid = io_input_valid_913; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_913_io_iormac = io_iormac_913; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_914_clock = clock;
  assign bc_pe_914_reset = reset;
  assign bc_pe_914_io_ho_input = bc_pe_913_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_914_io_ve_input = bc_pe_882_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_914_io_input_valid = io_input_valid_914; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_914_io_iormac = io_iormac_914; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_915_clock = clock;
  assign bc_pe_915_reset = reset;
  assign bc_pe_915_io_ho_input = bc_pe_914_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_915_io_ve_input = bc_pe_883_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_915_io_input_valid = io_input_valid_915; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_915_io_iormac = io_iormac_915; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_916_clock = clock;
  assign bc_pe_916_reset = reset;
  assign bc_pe_916_io_ho_input = bc_pe_915_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_916_io_ve_input = bc_pe_884_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_916_io_input_valid = io_input_valid_916; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_916_io_iormac = io_iormac_916; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_917_clock = clock;
  assign bc_pe_917_reset = reset;
  assign bc_pe_917_io_ho_input = bc_pe_916_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_917_io_ve_input = bc_pe_885_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_917_io_input_valid = io_input_valid_917; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_917_io_iormac = io_iormac_917; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_918_clock = clock;
  assign bc_pe_918_reset = reset;
  assign bc_pe_918_io_ho_input = bc_pe_917_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_918_io_ve_input = bc_pe_886_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_918_io_input_valid = io_input_valid_918; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_918_io_iormac = io_iormac_918; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_919_clock = clock;
  assign bc_pe_919_reset = reset;
  assign bc_pe_919_io_ho_input = bc_pe_918_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_919_io_ve_input = bc_pe_887_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_919_io_input_valid = io_input_valid_919; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_919_io_iormac = io_iormac_919; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_920_clock = clock;
  assign bc_pe_920_reset = reset;
  assign bc_pe_920_io_ho_input = bc_pe_919_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_920_io_ve_input = bc_pe_888_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_920_io_input_valid = io_input_valid_920; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_920_io_iormac = io_iormac_920; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_921_clock = clock;
  assign bc_pe_921_reset = reset;
  assign bc_pe_921_io_ho_input = bc_pe_920_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_921_io_ve_input = bc_pe_889_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_921_io_input_valid = io_input_valid_921; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_921_io_iormac = io_iormac_921; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_922_clock = clock;
  assign bc_pe_922_reset = reset;
  assign bc_pe_922_io_ho_input = bc_pe_921_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_922_io_ve_input = bc_pe_890_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_922_io_input_valid = io_input_valid_922; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_922_io_iormac = io_iormac_922; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_923_clock = clock;
  assign bc_pe_923_reset = reset;
  assign bc_pe_923_io_ho_input = bc_pe_922_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_923_io_ve_input = bc_pe_891_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_923_io_input_valid = io_input_valid_923; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_923_io_iormac = io_iormac_923; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_924_clock = clock;
  assign bc_pe_924_reset = reset;
  assign bc_pe_924_io_ho_input = bc_pe_923_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_924_io_ve_input = bc_pe_892_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_924_io_input_valid = io_input_valid_924; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_924_io_iormac = io_iormac_924; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_925_clock = clock;
  assign bc_pe_925_reset = reset;
  assign bc_pe_925_io_ho_input = bc_pe_924_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_925_io_ve_input = bc_pe_893_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_925_io_input_valid = io_input_valid_925; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_925_io_iormac = io_iormac_925; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_926_clock = clock;
  assign bc_pe_926_reset = reset;
  assign bc_pe_926_io_ho_input = bc_pe_925_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_926_io_ve_input = bc_pe_894_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_926_io_input_valid = io_input_valid_926; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_926_io_iormac = io_iormac_926; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_927_clock = clock;
  assign bc_pe_927_reset = reset;
  assign bc_pe_927_io_ho_input = bc_pe_926_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_927_io_ve_input = bc_pe_895_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_927_io_input_valid = io_input_valid_927; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_927_io_iormac = io_iormac_927; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_928_clock = clock;
  assign bc_pe_928_reset = reset;
  assign bc_pe_928_io_ho_input = io_x_input_29; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_928_io_ve_input = bc_pe_896_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_928_io_input_valid = io_input_valid_928; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_928_io_iormac = io_iormac_928; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_929_clock = clock;
  assign bc_pe_929_reset = reset;
  assign bc_pe_929_io_ho_input = bc_pe_928_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_929_io_ve_input = bc_pe_897_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_929_io_input_valid = io_input_valid_929; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_929_io_iormac = io_iormac_929; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_930_clock = clock;
  assign bc_pe_930_reset = reset;
  assign bc_pe_930_io_ho_input = bc_pe_929_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_930_io_ve_input = bc_pe_898_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_930_io_input_valid = io_input_valid_930; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_930_io_iormac = io_iormac_930; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_931_clock = clock;
  assign bc_pe_931_reset = reset;
  assign bc_pe_931_io_ho_input = bc_pe_930_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_931_io_ve_input = bc_pe_899_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_931_io_input_valid = io_input_valid_931; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_931_io_iormac = io_iormac_931; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_932_clock = clock;
  assign bc_pe_932_reset = reset;
  assign bc_pe_932_io_ho_input = bc_pe_931_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_932_io_ve_input = bc_pe_900_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_932_io_input_valid = io_input_valid_932; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_932_io_iormac = io_iormac_932; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_933_clock = clock;
  assign bc_pe_933_reset = reset;
  assign bc_pe_933_io_ho_input = bc_pe_932_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_933_io_ve_input = bc_pe_901_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_933_io_input_valid = io_input_valid_933; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_933_io_iormac = io_iormac_933; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_934_clock = clock;
  assign bc_pe_934_reset = reset;
  assign bc_pe_934_io_ho_input = bc_pe_933_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_934_io_ve_input = bc_pe_902_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_934_io_input_valid = io_input_valid_934; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_934_io_iormac = io_iormac_934; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_935_clock = clock;
  assign bc_pe_935_reset = reset;
  assign bc_pe_935_io_ho_input = bc_pe_934_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_935_io_ve_input = bc_pe_903_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_935_io_input_valid = io_input_valid_935; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_935_io_iormac = io_iormac_935; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_936_clock = clock;
  assign bc_pe_936_reset = reset;
  assign bc_pe_936_io_ho_input = bc_pe_935_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_936_io_ve_input = bc_pe_904_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_936_io_input_valid = io_input_valid_936; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_936_io_iormac = io_iormac_936; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_937_clock = clock;
  assign bc_pe_937_reset = reset;
  assign bc_pe_937_io_ho_input = bc_pe_936_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_937_io_ve_input = bc_pe_905_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_937_io_input_valid = io_input_valid_937; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_937_io_iormac = io_iormac_937; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_938_clock = clock;
  assign bc_pe_938_reset = reset;
  assign bc_pe_938_io_ho_input = bc_pe_937_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_938_io_ve_input = bc_pe_906_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_938_io_input_valid = io_input_valid_938; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_938_io_iormac = io_iormac_938; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_939_clock = clock;
  assign bc_pe_939_reset = reset;
  assign bc_pe_939_io_ho_input = bc_pe_938_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_939_io_ve_input = bc_pe_907_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_939_io_input_valid = io_input_valid_939; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_939_io_iormac = io_iormac_939; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_940_clock = clock;
  assign bc_pe_940_reset = reset;
  assign bc_pe_940_io_ho_input = bc_pe_939_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_940_io_ve_input = bc_pe_908_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_940_io_input_valid = io_input_valid_940; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_940_io_iormac = io_iormac_940; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_941_clock = clock;
  assign bc_pe_941_reset = reset;
  assign bc_pe_941_io_ho_input = bc_pe_940_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_941_io_ve_input = bc_pe_909_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_941_io_input_valid = io_input_valid_941; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_941_io_iormac = io_iormac_941; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_942_clock = clock;
  assign bc_pe_942_reset = reset;
  assign bc_pe_942_io_ho_input = bc_pe_941_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_942_io_ve_input = bc_pe_910_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_942_io_input_valid = io_input_valid_942; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_942_io_iormac = io_iormac_942; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_943_clock = clock;
  assign bc_pe_943_reset = reset;
  assign bc_pe_943_io_ho_input = bc_pe_942_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_943_io_ve_input = bc_pe_911_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_943_io_input_valid = io_input_valid_943; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_943_io_iormac = io_iormac_943; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_944_clock = clock;
  assign bc_pe_944_reset = reset;
  assign bc_pe_944_io_ho_input = bc_pe_943_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_944_io_ve_input = bc_pe_912_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_944_io_input_valid = io_input_valid_944; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_944_io_iormac = io_iormac_944; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_945_clock = clock;
  assign bc_pe_945_reset = reset;
  assign bc_pe_945_io_ho_input = bc_pe_944_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_945_io_ve_input = bc_pe_913_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_945_io_input_valid = io_input_valid_945; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_945_io_iormac = io_iormac_945; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_946_clock = clock;
  assign bc_pe_946_reset = reset;
  assign bc_pe_946_io_ho_input = bc_pe_945_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_946_io_ve_input = bc_pe_914_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_946_io_input_valid = io_input_valid_946; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_946_io_iormac = io_iormac_946; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_947_clock = clock;
  assign bc_pe_947_reset = reset;
  assign bc_pe_947_io_ho_input = bc_pe_946_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_947_io_ve_input = bc_pe_915_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_947_io_input_valid = io_input_valid_947; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_947_io_iormac = io_iormac_947; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_948_clock = clock;
  assign bc_pe_948_reset = reset;
  assign bc_pe_948_io_ho_input = bc_pe_947_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_948_io_ve_input = bc_pe_916_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_948_io_input_valid = io_input_valid_948; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_948_io_iormac = io_iormac_948; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_949_clock = clock;
  assign bc_pe_949_reset = reset;
  assign bc_pe_949_io_ho_input = bc_pe_948_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_949_io_ve_input = bc_pe_917_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_949_io_input_valid = io_input_valid_949; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_949_io_iormac = io_iormac_949; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_950_clock = clock;
  assign bc_pe_950_reset = reset;
  assign bc_pe_950_io_ho_input = bc_pe_949_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_950_io_ve_input = bc_pe_918_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_950_io_input_valid = io_input_valid_950; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_950_io_iormac = io_iormac_950; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_951_clock = clock;
  assign bc_pe_951_reset = reset;
  assign bc_pe_951_io_ho_input = bc_pe_950_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_951_io_ve_input = bc_pe_919_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_951_io_input_valid = io_input_valid_951; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_951_io_iormac = io_iormac_951; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_952_clock = clock;
  assign bc_pe_952_reset = reset;
  assign bc_pe_952_io_ho_input = bc_pe_951_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_952_io_ve_input = bc_pe_920_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_952_io_input_valid = io_input_valid_952; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_952_io_iormac = io_iormac_952; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_953_clock = clock;
  assign bc_pe_953_reset = reset;
  assign bc_pe_953_io_ho_input = bc_pe_952_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_953_io_ve_input = bc_pe_921_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_953_io_input_valid = io_input_valid_953; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_953_io_iormac = io_iormac_953; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_954_clock = clock;
  assign bc_pe_954_reset = reset;
  assign bc_pe_954_io_ho_input = bc_pe_953_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_954_io_ve_input = bc_pe_922_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_954_io_input_valid = io_input_valid_954; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_954_io_iormac = io_iormac_954; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_955_clock = clock;
  assign bc_pe_955_reset = reset;
  assign bc_pe_955_io_ho_input = bc_pe_954_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_955_io_ve_input = bc_pe_923_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_955_io_input_valid = io_input_valid_955; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_955_io_iormac = io_iormac_955; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_956_clock = clock;
  assign bc_pe_956_reset = reset;
  assign bc_pe_956_io_ho_input = bc_pe_955_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_956_io_ve_input = bc_pe_924_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_956_io_input_valid = io_input_valid_956; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_956_io_iormac = io_iormac_956; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_957_clock = clock;
  assign bc_pe_957_reset = reset;
  assign bc_pe_957_io_ho_input = bc_pe_956_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_957_io_ve_input = bc_pe_925_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_957_io_input_valid = io_input_valid_957; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_957_io_iormac = io_iormac_957; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_958_clock = clock;
  assign bc_pe_958_reset = reset;
  assign bc_pe_958_io_ho_input = bc_pe_957_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_958_io_ve_input = bc_pe_926_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_958_io_input_valid = io_input_valid_958; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_958_io_iormac = io_iormac_958; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_959_clock = clock;
  assign bc_pe_959_reset = reset;
  assign bc_pe_959_io_ho_input = bc_pe_958_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_959_io_ve_input = bc_pe_927_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_959_io_input_valid = io_input_valid_959; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_959_io_iormac = io_iormac_959; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_960_clock = clock;
  assign bc_pe_960_reset = reset;
  assign bc_pe_960_io_ho_input = io_x_input_30; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_960_io_ve_input = bc_pe_928_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_960_io_input_valid = io_input_valid_960; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_960_io_iormac = io_iormac_960; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_961_clock = clock;
  assign bc_pe_961_reset = reset;
  assign bc_pe_961_io_ho_input = bc_pe_960_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_961_io_ve_input = bc_pe_929_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_961_io_input_valid = io_input_valid_961; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_961_io_iormac = io_iormac_961; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_962_clock = clock;
  assign bc_pe_962_reset = reset;
  assign bc_pe_962_io_ho_input = bc_pe_961_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_962_io_ve_input = bc_pe_930_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_962_io_input_valid = io_input_valid_962; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_962_io_iormac = io_iormac_962; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_963_clock = clock;
  assign bc_pe_963_reset = reset;
  assign bc_pe_963_io_ho_input = bc_pe_962_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_963_io_ve_input = bc_pe_931_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_963_io_input_valid = io_input_valid_963; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_963_io_iormac = io_iormac_963; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_964_clock = clock;
  assign bc_pe_964_reset = reset;
  assign bc_pe_964_io_ho_input = bc_pe_963_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_964_io_ve_input = bc_pe_932_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_964_io_input_valid = io_input_valid_964; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_964_io_iormac = io_iormac_964; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_965_clock = clock;
  assign bc_pe_965_reset = reset;
  assign bc_pe_965_io_ho_input = bc_pe_964_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_965_io_ve_input = bc_pe_933_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_965_io_input_valid = io_input_valid_965; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_965_io_iormac = io_iormac_965; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_966_clock = clock;
  assign bc_pe_966_reset = reset;
  assign bc_pe_966_io_ho_input = bc_pe_965_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_966_io_ve_input = bc_pe_934_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_966_io_input_valid = io_input_valid_966; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_966_io_iormac = io_iormac_966; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_967_clock = clock;
  assign bc_pe_967_reset = reset;
  assign bc_pe_967_io_ho_input = bc_pe_966_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_967_io_ve_input = bc_pe_935_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_967_io_input_valid = io_input_valid_967; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_967_io_iormac = io_iormac_967; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_968_clock = clock;
  assign bc_pe_968_reset = reset;
  assign bc_pe_968_io_ho_input = bc_pe_967_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_968_io_ve_input = bc_pe_936_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_968_io_input_valid = io_input_valid_968; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_968_io_iormac = io_iormac_968; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_969_clock = clock;
  assign bc_pe_969_reset = reset;
  assign bc_pe_969_io_ho_input = bc_pe_968_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_969_io_ve_input = bc_pe_937_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_969_io_input_valid = io_input_valid_969; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_969_io_iormac = io_iormac_969; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_970_clock = clock;
  assign bc_pe_970_reset = reset;
  assign bc_pe_970_io_ho_input = bc_pe_969_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_970_io_ve_input = bc_pe_938_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_970_io_input_valid = io_input_valid_970; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_970_io_iormac = io_iormac_970; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_971_clock = clock;
  assign bc_pe_971_reset = reset;
  assign bc_pe_971_io_ho_input = bc_pe_970_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_971_io_ve_input = bc_pe_939_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_971_io_input_valid = io_input_valid_971; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_971_io_iormac = io_iormac_971; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_972_clock = clock;
  assign bc_pe_972_reset = reset;
  assign bc_pe_972_io_ho_input = bc_pe_971_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_972_io_ve_input = bc_pe_940_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_972_io_input_valid = io_input_valid_972; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_972_io_iormac = io_iormac_972; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_973_clock = clock;
  assign bc_pe_973_reset = reset;
  assign bc_pe_973_io_ho_input = bc_pe_972_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_973_io_ve_input = bc_pe_941_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_973_io_input_valid = io_input_valid_973; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_973_io_iormac = io_iormac_973; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_974_clock = clock;
  assign bc_pe_974_reset = reset;
  assign bc_pe_974_io_ho_input = bc_pe_973_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_974_io_ve_input = bc_pe_942_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_974_io_input_valid = io_input_valid_974; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_974_io_iormac = io_iormac_974; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_975_clock = clock;
  assign bc_pe_975_reset = reset;
  assign bc_pe_975_io_ho_input = bc_pe_974_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_975_io_ve_input = bc_pe_943_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_975_io_input_valid = io_input_valid_975; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_975_io_iormac = io_iormac_975; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_976_clock = clock;
  assign bc_pe_976_reset = reset;
  assign bc_pe_976_io_ho_input = bc_pe_975_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_976_io_ve_input = bc_pe_944_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_976_io_input_valid = io_input_valid_976; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_976_io_iormac = io_iormac_976; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_977_clock = clock;
  assign bc_pe_977_reset = reset;
  assign bc_pe_977_io_ho_input = bc_pe_976_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_977_io_ve_input = bc_pe_945_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_977_io_input_valid = io_input_valid_977; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_977_io_iormac = io_iormac_977; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_978_clock = clock;
  assign bc_pe_978_reset = reset;
  assign bc_pe_978_io_ho_input = bc_pe_977_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_978_io_ve_input = bc_pe_946_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_978_io_input_valid = io_input_valid_978; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_978_io_iormac = io_iormac_978; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_979_clock = clock;
  assign bc_pe_979_reset = reset;
  assign bc_pe_979_io_ho_input = bc_pe_978_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_979_io_ve_input = bc_pe_947_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_979_io_input_valid = io_input_valid_979; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_979_io_iormac = io_iormac_979; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_980_clock = clock;
  assign bc_pe_980_reset = reset;
  assign bc_pe_980_io_ho_input = bc_pe_979_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_980_io_ve_input = bc_pe_948_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_980_io_input_valid = io_input_valid_980; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_980_io_iormac = io_iormac_980; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_981_clock = clock;
  assign bc_pe_981_reset = reset;
  assign bc_pe_981_io_ho_input = bc_pe_980_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_981_io_ve_input = bc_pe_949_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_981_io_input_valid = io_input_valid_981; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_981_io_iormac = io_iormac_981; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_982_clock = clock;
  assign bc_pe_982_reset = reset;
  assign bc_pe_982_io_ho_input = bc_pe_981_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_982_io_ve_input = bc_pe_950_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_982_io_input_valid = io_input_valid_982; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_982_io_iormac = io_iormac_982; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_983_clock = clock;
  assign bc_pe_983_reset = reset;
  assign bc_pe_983_io_ho_input = bc_pe_982_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_983_io_ve_input = bc_pe_951_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_983_io_input_valid = io_input_valid_983; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_983_io_iormac = io_iormac_983; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_984_clock = clock;
  assign bc_pe_984_reset = reset;
  assign bc_pe_984_io_ho_input = bc_pe_983_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_984_io_ve_input = bc_pe_952_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_984_io_input_valid = io_input_valid_984; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_984_io_iormac = io_iormac_984; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_985_clock = clock;
  assign bc_pe_985_reset = reset;
  assign bc_pe_985_io_ho_input = bc_pe_984_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_985_io_ve_input = bc_pe_953_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_985_io_input_valid = io_input_valid_985; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_985_io_iormac = io_iormac_985; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_986_clock = clock;
  assign bc_pe_986_reset = reset;
  assign bc_pe_986_io_ho_input = bc_pe_985_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_986_io_ve_input = bc_pe_954_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_986_io_input_valid = io_input_valid_986; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_986_io_iormac = io_iormac_986; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_987_clock = clock;
  assign bc_pe_987_reset = reset;
  assign bc_pe_987_io_ho_input = bc_pe_986_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_987_io_ve_input = bc_pe_955_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_987_io_input_valid = io_input_valid_987; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_987_io_iormac = io_iormac_987; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_988_clock = clock;
  assign bc_pe_988_reset = reset;
  assign bc_pe_988_io_ho_input = bc_pe_987_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_988_io_ve_input = bc_pe_956_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_988_io_input_valid = io_input_valid_988; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_988_io_iormac = io_iormac_988; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_989_clock = clock;
  assign bc_pe_989_reset = reset;
  assign bc_pe_989_io_ho_input = bc_pe_988_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_989_io_ve_input = bc_pe_957_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_989_io_input_valid = io_input_valid_989; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_989_io_iormac = io_iormac_989; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_990_clock = clock;
  assign bc_pe_990_reset = reset;
  assign bc_pe_990_io_ho_input = bc_pe_989_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_990_io_ve_input = bc_pe_958_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_990_io_input_valid = io_input_valid_990; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_990_io_iormac = io_iormac_990; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_991_clock = clock;
  assign bc_pe_991_reset = reset;
  assign bc_pe_991_io_ho_input = bc_pe_990_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_991_io_ve_input = bc_pe_959_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_991_io_input_valid = io_input_valid_991; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_991_io_iormac = io_iormac_991; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_992_clock = clock;
  assign bc_pe_992_reset = reset;
  assign bc_pe_992_io_ho_input = io_x_input_31; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_992_io_ve_input = bc_pe_960_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_992_io_input_valid = io_input_valid_992; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_992_io_iormac = io_iormac_992; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_993_clock = clock;
  assign bc_pe_993_reset = reset;
  assign bc_pe_993_io_ho_input = bc_pe_992_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_993_io_ve_input = bc_pe_961_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_993_io_input_valid = io_input_valid_993; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_993_io_iormac = io_iormac_993; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_994_clock = clock;
  assign bc_pe_994_reset = reset;
  assign bc_pe_994_io_ho_input = bc_pe_993_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_994_io_ve_input = bc_pe_962_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_994_io_input_valid = io_input_valid_994; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_994_io_iormac = io_iormac_994; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_995_clock = clock;
  assign bc_pe_995_reset = reset;
  assign bc_pe_995_io_ho_input = bc_pe_994_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_995_io_ve_input = bc_pe_963_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_995_io_input_valid = io_input_valid_995; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_995_io_iormac = io_iormac_995; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_996_clock = clock;
  assign bc_pe_996_reset = reset;
  assign bc_pe_996_io_ho_input = bc_pe_995_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_996_io_ve_input = bc_pe_964_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_996_io_input_valid = io_input_valid_996; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_996_io_iormac = io_iormac_996; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_997_clock = clock;
  assign bc_pe_997_reset = reset;
  assign bc_pe_997_io_ho_input = bc_pe_996_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_997_io_ve_input = bc_pe_965_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_997_io_input_valid = io_input_valid_997; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_997_io_iormac = io_iormac_997; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_998_clock = clock;
  assign bc_pe_998_reset = reset;
  assign bc_pe_998_io_ho_input = bc_pe_997_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_998_io_ve_input = bc_pe_966_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_998_io_input_valid = io_input_valid_998; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_998_io_iormac = io_iormac_998; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_999_clock = clock;
  assign bc_pe_999_reset = reset;
  assign bc_pe_999_io_ho_input = bc_pe_998_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_999_io_ve_input = bc_pe_967_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_999_io_input_valid = io_input_valid_999; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_999_io_iormac = io_iormac_999; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1000_clock = clock;
  assign bc_pe_1000_reset = reset;
  assign bc_pe_1000_io_ho_input = bc_pe_999_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1000_io_ve_input = bc_pe_968_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1000_io_input_valid = io_input_valid_1000; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1000_io_iormac = io_iormac_1000; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1001_clock = clock;
  assign bc_pe_1001_reset = reset;
  assign bc_pe_1001_io_ho_input = bc_pe_1000_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1001_io_ve_input = bc_pe_969_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1001_io_input_valid = io_input_valid_1001; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1001_io_iormac = io_iormac_1001; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1002_clock = clock;
  assign bc_pe_1002_reset = reset;
  assign bc_pe_1002_io_ho_input = bc_pe_1001_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1002_io_ve_input = bc_pe_970_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1002_io_input_valid = io_input_valid_1002; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1002_io_iormac = io_iormac_1002; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1003_clock = clock;
  assign bc_pe_1003_reset = reset;
  assign bc_pe_1003_io_ho_input = bc_pe_1002_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1003_io_ve_input = bc_pe_971_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1003_io_input_valid = io_input_valid_1003; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1003_io_iormac = io_iormac_1003; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1004_clock = clock;
  assign bc_pe_1004_reset = reset;
  assign bc_pe_1004_io_ho_input = bc_pe_1003_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1004_io_ve_input = bc_pe_972_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1004_io_input_valid = io_input_valid_1004; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1004_io_iormac = io_iormac_1004; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1005_clock = clock;
  assign bc_pe_1005_reset = reset;
  assign bc_pe_1005_io_ho_input = bc_pe_1004_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1005_io_ve_input = bc_pe_973_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1005_io_input_valid = io_input_valid_1005; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1005_io_iormac = io_iormac_1005; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1006_clock = clock;
  assign bc_pe_1006_reset = reset;
  assign bc_pe_1006_io_ho_input = bc_pe_1005_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1006_io_ve_input = bc_pe_974_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1006_io_input_valid = io_input_valid_1006; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1006_io_iormac = io_iormac_1006; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1007_clock = clock;
  assign bc_pe_1007_reset = reset;
  assign bc_pe_1007_io_ho_input = bc_pe_1006_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1007_io_ve_input = bc_pe_975_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1007_io_input_valid = io_input_valid_1007; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1007_io_iormac = io_iormac_1007; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1008_clock = clock;
  assign bc_pe_1008_reset = reset;
  assign bc_pe_1008_io_ho_input = bc_pe_1007_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1008_io_ve_input = bc_pe_976_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1008_io_input_valid = io_input_valid_1008; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1008_io_iormac = io_iormac_1008; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1009_clock = clock;
  assign bc_pe_1009_reset = reset;
  assign bc_pe_1009_io_ho_input = bc_pe_1008_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1009_io_ve_input = bc_pe_977_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1009_io_input_valid = io_input_valid_1009; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1009_io_iormac = io_iormac_1009; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1010_clock = clock;
  assign bc_pe_1010_reset = reset;
  assign bc_pe_1010_io_ho_input = bc_pe_1009_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1010_io_ve_input = bc_pe_978_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1010_io_input_valid = io_input_valid_1010; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1010_io_iormac = io_iormac_1010; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1011_clock = clock;
  assign bc_pe_1011_reset = reset;
  assign bc_pe_1011_io_ho_input = bc_pe_1010_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1011_io_ve_input = bc_pe_979_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1011_io_input_valid = io_input_valid_1011; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1011_io_iormac = io_iormac_1011; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1012_clock = clock;
  assign bc_pe_1012_reset = reset;
  assign bc_pe_1012_io_ho_input = bc_pe_1011_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1012_io_ve_input = bc_pe_980_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1012_io_input_valid = io_input_valid_1012; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1012_io_iormac = io_iormac_1012; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1013_clock = clock;
  assign bc_pe_1013_reset = reset;
  assign bc_pe_1013_io_ho_input = bc_pe_1012_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1013_io_ve_input = bc_pe_981_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1013_io_input_valid = io_input_valid_1013; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1013_io_iormac = io_iormac_1013; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1014_clock = clock;
  assign bc_pe_1014_reset = reset;
  assign bc_pe_1014_io_ho_input = bc_pe_1013_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1014_io_ve_input = bc_pe_982_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1014_io_input_valid = io_input_valid_1014; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1014_io_iormac = io_iormac_1014; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1015_clock = clock;
  assign bc_pe_1015_reset = reset;
  assign bc_pe_1015_io_ho_input = bc_pe_1014_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1015_io_ve_input = bc_pe_983_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1015_io_input_valid = io_input_valid_1015; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1015_io_iormac = io_iormac_1015; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1016_clock = clock;
  assign bc_pe_1016_reset = reset;
  assign bc_pe_1016_io_ho_input = bc_pe_1015_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1016_io_ve_input = bc_pe_984_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1016_io_input_valid = io_input_valid_1016; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1016_io_iormac = io_iormac_1016; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1017_clock = clock;
  assign bc_pe_1017_reset = reset;
  assign bc_pe_1017_io_ho_input = bc_pe_1016_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1017_io_ve_input = bc_pe_985_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1017_io_input_valid = io_input_valid_1017; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1017_io_iormac = io_iormac_1017; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1018_clock = clock;
  assign bc_pe_1018_reset = reset;
  assign bc_pe_1018_io_ho_input = bc_pe_1017_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1018_io_ve_input = bc_pe_986_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1018_io_input_valid = io_input_valid_1018; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1018_io_iormac = io_iormac_1018; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1019_clock = clock;
  assign bc_pe_1019_reset = reset;
  assign bc_pe_1019_io_ho_input = bc_pe_1018_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1019_io_ve_input = bc_pe_987_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1019_io_input_valid = io_input_valid_1019; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1019_io_iormac = io_iormac_1019; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1020_clock = clock;
  assign bc_pe_1020_reset = reset;
  assign bc_pe_1020_io_ho_input = bc_pe_1019_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1020_io_ve_input = bc_pe_988_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1020_io_input_valid = io_input_valid_1020; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1020_io_iormac = io_iormac_1020; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1021_clock = clock;
  assign bc_pe_1021_reset = reset;
  assign bc_pe_1021_io_ho_input = bc_pe_1020_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1021_io_ve_input = bc_pe_989_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1021_io_input_valid = io_input_valid_1021; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1021_io_iormac = io_iormac_1021; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1022_clock = clock;
  assign bc_pe_1022_reset = reset;
  assign bc_pe_1022_io_ho_input = bc_pe_1021_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1022_io_ve_input = bc_pe_990_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1022_io_input_valid = io_input_valid_1022; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1022_io_iormac = io_iormac_1022; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_1023_clock = clock;
  assign bc_pe_1023_reset = reset;
  assign bc_pe_1023_io_ho_input = bc_pe_1022_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1023_io_ve_input = bc_pe_991_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1023_io_input_valid = io_input_valid_1023; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_1023_io_iormac = io_iormac_1023; // @[bc_mmul.scala 22:28 78:47]
endmodule
