module bc_pe(
  input         clock,
  input         reset,
  input  [15:0] io_ho_input,
  input  [31:0] io_ve_input,
  input         io_input_valid,
  input         io_iormac,
  output [31:0] io_ve_out,
  output [15:0] io_ho_out,
  output [31:0] io_res_out
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] mac; // @[bc_pe.scala 30:23]
  reg [15:0] ho_reg; // @[bc_pe.scala 31:23]
  reg [31:0] ve_reg; // @[bc_pe.scala 32:23]
  reg  REG; // @[bc_pe.scala 37:42]
  wire  _T_1 = io_input_valid & ~REG; // @[bc_pe.scala 37:31]
  wire [47:0] _mac_T = io_ho_input * io_ve_input; // @[bc_pe.scala 44:39]
  wire [47:0] _GEN_3 = {{16'd0}, mac}; // @[bc_pe.scala 44:24]
  wire [47:0] _mac_T_2 = _GEN_3 + _mac_T; // @[bc_pe.scala 44:24]
  wire [47:0] _GEN_0 = _T_1 ? _mac_T_2 : {{16'd0}, mac}; // @[bc_pe.scala 42:46 44:17 30:23]
  wire [47:0] _GEN_4 = reset ? 48'h0 : _GEN_0; // @[bc_pe.scala 30:{23,23}]
  assign io_ve_out = io_iormac ? ve_reg : mac; // @[bc_pe.scala 51:20]
  assign io_ho_out = ho_reg; // @[bc_pe.scala 52:14]
  assign io_res_out = mac; // @[bc_pe.scala 50:14]
  always @(posedge clock) begin
    mac <= _GEN_4[31:0]; // @[bc_pe.scala 30:{23,23}]
    if (reset) begin // @[bc_pe.scala 31:23]
      ho_reg <= 16'h0; // @[bc_pe.scala 31:23]
    end else if (_T_1) begin // @[bc_pe.scala 42:46]
      ho_reg <= io_ho_input; // @[bc_pe.scala 45:17]
    end
    if (reset) begin // @[bc_pe.scala 32:23]
      ve_reg <= 32'h0; // @[bc_pe.scala 32:23]
    end else if (_T_1) begin // @[bc_pe.scala 42:46]
      ve_reg <= io_ve_input; // @[bc_pe.scala 46:17]
    end
    REG <= io_input_valid; // @[bc_pe.scala 37:42]
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  mac = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  ho_reg = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  ve_reg = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  REG = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module bc_mmul(
  input         clock,
  input         reset,
  input  [15:0] io_x_input_0,
  input  [15:0] io_x_input_1,
  input  [15:0] io_x_input_2,
  input  [15:0] io_x_input_3,
  input  [15:0] io_x_input_4,
  input  [15:0] io_x_input_5,
  input  [15:0] io_x_input_6,
  input  [15:0] io_x_input_7,
  input  [15:0] io_x_input_8,
  input  [15:0] io_x_input_9,
  input  [15:0] io_x_input_10,
  input  [15:0] io_x_input_11,
  input  [15:0] io_x_input_12,
  input  [15:0] io_x_input_13,
  input  [15:0] io_x_input_14,
  input  [15:0] io_x_input_15,
  input  [31:0] io_w_input_0,
  input  [31:0] io_w_input_1,
  input  [31:0] io_w_input_2,
  input  [31:0] io_w_input_3,
  input  [31:0] io_w_input_4,
  input  [31:0] io_w_input_5,
  input  [31:0] io_w_input_6,
  input  [31:0] io_w_input_7,
  input  [31:0] io_w_input_8,
  input  [31:0] io_w_input_9,
  input  [31:0] io_w_input_10,
  input  [31:0] io_w_input_11,
  input  [31:0] io_w_input_12,
  input  [31:0] io_w_input_13,
  input  [31:0] io_w_input_14,
  input  [31:0] io_w_input_15,
  input         io_input_valid_0,
  input         io_input_valid_1,
  input         io_input_valid_2,
  input         io_input_valid_3,
  input         io_input_valid_4,
  input         io_input_valid_5,
  input         io_input_valid_6,
  input         io_input_valid_7,
  input         io_input_valid_8,
  input         io_input_valid_9,
  input         io_input_valid_10,
  input         io_input_valid_11,
  input         io_input_valid_12,
  input         io_input_valid_13,
  input         io_input_valid_14,
  input         io_input_valid_15,
  input         io_input_valid_16,
  input         io_input_valid_17,
  input         io_input_valid_18,
  input         io_input_valid_19,
  input         io_input_valid_20,
  input         io_input_valid_21,
  input         io_input_valid_22,
  input         io_input_valid_23,
  input         io_input_valid_24,
  input         io_input_valid_25,
  input         io_input_valid_26,
  input         io_input_valid_27,
  input         io_input_valid_28,
  input         io_input_valid_29,
  input         io_input_valid_30,
  input         io_input_valid_31,
  input         io_input_valid_32,
  input         io_input_valid_33,
  input         io_input_valid_34,
  input         io_input_valid_35,
  input         io_input_valid_36,
  input         io_input_valid_37,
  input         io_input_valid_38,
  input         io_input_valid_39,
  input         io_input_valid_40,
  input         io_input_valid_41,
  input         io_input_valid_42,
  input         io_input_valid_43,
  input         io_input_valid_44,
  input         io_input_valid_45,
  input         io_input_valid_46,
  input         io_input_valid_47,
  input         io_input_valid_48,
  input         io_input_valid_49,
  input         io_input_valid_50,
  input         io_input_valid_51,
  input         io_input_valid_52,
  input         io_input_valid_53,
  input         io_input_valid_54,
  input         io_input_valid_55,
  input         io_input_valid_56,
  input         io_input_valid_57,
  input         io_input_valid_58,
  input         io_input_valid_59,
  input         io_input_valid_60,
  input         io_input_valid_61,
  input         io_input_valid_62,
  input         io_input_valid_63,
  input         io_input_valid_64,
  input         io_input_valid_65,
  input         io_input_valid_66,
  input         io_input_valid_67,
  input         io_input_valid_68,
  input         io_input_valid_69,
  input         io_input_valid_70,
  input         io_input_valid_71,
  input         io_input_valid_72,
  input         io_input_valid_73,
  input         io_input_valid_74,
  input         io_input_valid_75,
  input         io_input_valid_76,
  input         io_input_valid_77,
  input         io_input_valid_78,
  input         io_input_valid_79,
  input         io_input_valid_80,
  input         io_input_valid_81,
  input         io_input_valid_82,
  input         io_input_valid_83,
  input         io_input_valid_84,
  input         io_input_valid_85,
  input         io_input_valid_86,
  input         io_input_valid_87,
  input         io_input_valid_88,
  input         io_input_valid_89,
  input         io_input_valid_90,
  input         io_input_valid_91,
  input         io_input_valid_92,
  input         io_input_valid_93,
  input         io_input_valid_94,
  input         io_input_valid_95,
  input         io_input_valid_96,
  input         io_input_valid_97,
  input         io_input_valid_98,
  input         io_input_valid_99,
  input         io_input_valid_100,
  input         io_input_valid_101,
  input         io_input_valid_102,
  input         io_input_valid_103,
  input         io_input_valid_104,
  input         io_input_valid_105,
  input         io_input_valid_106,
  input         io_input_valid_107,
  input         io_input_valid_108,
  input         io_input_valid_109,
  input         io_input_valid_110,
  input         io_input_valid_111,
  input         io_input_valid_112,
  input         io_input_valid_113,
  input         io_input_valid_114,
  input         io_input_valid_115,
  input         io_input_valid_116,
  input         io_input_valid_117,
  input         io_input_valid_118,
  input         io_input_valid_119,
  input         io_input_valid_120,
  input         io_input_valid_121,
  input         io_input_valid_122,
  input         io_input_valid_123,
  input         io_input_valid_124,
  input         io_input_valid_125,
  input         io_input_valid_126,
  input         io_input_valid_127,
  input         io_input_valid_128,
  input         io_input_valid_129,
  input         io_input_valid_130,
  input         io_input_valid_131,
  input         io_input_valid_132,
  input         io_input_valid_133,
  input         io_input_valid_134,
  input         io_input_valid_135,
  input         io_input_valid_136,
  input         io_input_valid_137,
  input         io_input_valid_138,
  input         io_input_valid_139,
  input         io_input_valid_140,
  input         io_input_valid_141,
  input         io_input_valid_142,
  input         io_input_valid_143,
  input         io_input_valid_144,
  input         io_input_valid_145,
  input         io_input_valid_146,
  input         io_input_valid_147,
  input         io_input_valid_148,
  input         io_input_valid_149,
  input         io_input_valid_150,
  input         io_input_valid_151,
  input         io_input_valid_152,
  input         io_input_valid_153,
  input         io_input_valid_154,
  input         io_input_valid_155,
  input         io_input_valid_156,
  input         io_input_valid_157,
  input         io_input_valid_158,
  input         io_input_valid_159,
  input         io_input_valid_160,
  input         io_input_valid_161,
  input         io_input_valid_162,
  input         io_input_valid_163,
  input         io_input_valid_164,
  input         io_input_valid_165,
  input         io_input_valid_166,
  input         io_input_valid_167,
  input         io_input_valid_168,
  input         io_input_valid_169,
  input         io_input_valid_170,
  input         io_input_valid_171,
  input         io_input_valid_172,
  input         io_input_valid_173,
  input         io_input_valid_174,
  input         io_input_valid_175,
  input         io_input_valid_176,
  input         io_input_valid_177,
  input         io_input_valid_178,
  input         io_input_valid_179,
  input         io_input_valid_180,
  input         io_input_valid_181,
  input         io_input_valid_182,
  input         io_input_valid_183,
  input         io_input_valid_184,
  input         io_input_valid_185,
  input         io_input_valid_186,
  input         io_input_valid_187,
  input         io_input_valid_188,
  input         io_input_valid_189,
  input         io_input_valid_190,
  input         io_input_valid_191,
  input         io_input_valid_192,
  input         io_input_valid_193,
  input         io_input_valid_194,
  input         io_input_valid_195,
  input         io_input_valid_196,
  input         io_input_valid_197,
  input         io_input_valid_198,
  input         io_input_valid_199,
  input         io_input_valid_200,
  input         io_input_valid_201,
  input         io_input_valid_202,
  input         io_input_valid_203,
  input         io_input_valid_204,
  input         io_input_valid_205,
  input         io_input_valid_206,
  input         io_input_valid_207,
  input         io_input_valid_208,
  input         io_input_valid_209,
  input         io_input_valid_210,
  input         io_input_valid_211,
  input         io_input_valid_212,
  input         io_input_valid_213,
  input         io_input_valid_214,
  input         io_input_valid_215,
  input         io_input_valid_216,
  input         io_input_valid_217,
  input         io_input_valid_218,
  input         io_input_valid_219,
  input         io_input_valid_220,
  input         io_input_valid_221,
  input         io_input_valid_222,
  input         io_input_valid_223,
  input         io_input_valid_224,
  input         io_input_valid_225,
  input         io_input_valid_226,
  input         io_input_valid_227,
  input         io_input_valid_228,
  input         io_input_valid_229,
  input         io_input_valid_230,
  input         io_input_valid_231,
  input         io_input_valid_232,
  input         io_input_valid_233,
  input         io_input_valid_234,
  input         io_input_valid_235,
  input         io_input_valid_236,
  input         io_input_valid_237,
  input         io_input_valid_238,
  input         io_input_valid_239,
  input         io_input_valid_240,
  input         io_input_valid_241,
  input         io_input_valid_242,
  input         io_input_valid_243,
  input         io_input_valid_244,
  input         io_input_valid_245,
  input         io_input_valid_246,
  input         io_input_valid_247,
  input         io_input_valid_248,
  input         io_input_valid_249,
  input         io_input_valid_250,
  input         io_input_valid_251,
  input         io_input_valid_252,
  input         io_input_valid_253,
  input         io_input_valid_254,
  input         io_input_valid_255,
  input         io_iormac_0,
  input         io_iormac_1,
  input         io_iormac_2,
  input         io_iormac_3,
  input         io_iormac_4,
  input         io_iormac_5,
  input         io_iormac_6,
  input         io_iormac_7,
  input         io_iormac_8,
  input         io_iormac_9,
  input         io_iormac_10,
  input         io_iormac_11,
  input         io_iormac_12,
  input         io_iormac_13,
  input         io_iormac_14,
  input         io_iormac_15,
  input         io_iormac_16,
  input         io_iormac_17,
  input         io_iormac_18,
  input         io_iormac_19,
  input         io_iormac_20,
  input         io_iormac_21,
  input         io_iormac_22,
  input         io_iormac_23,
  input         io_iormac_24,
  input         io_iormac_25,
  input         io_iormac_26,
  input         io_iormac_27,
  input         io_iormac_28,
  input         io_iormac_29,
  input         io_iormac_30,
  input         io_iormac_31,
  input         io_iormac_32,
  input         io_iormac_33,
  input         io_iormac_34,
  input         io_iormac_35,
  input         io_iormac_36,
  input         io_iormac_37,
  input         io_iormac_38,
  input         io_iormac_39,
  input         io_iormac_40,
  input         io_iormac_41,
  input         io_iormac_42,
  input         io_iormac_43,
  input         io_iormac_44,
  input         io_iormac_45,
  input         io_iormac_46,
  input         io_iormac_47,
  input         io_iormac_48,
  input         io_iormac_49,
  input         io_iormac_50,
  input         io_iormac_51,
  input         io_iormac_52,
  input         io_iormac_53,
  input         io_iormac_54,
  input         io_iormac_55,
  input         io_iormac_56,
  input         io_iormac_57,
  input         io_iormac_58,
  input         io_iormac_59,
  input         io_iormac_60,
  input         io_iormac_61,
  input         io_iormac_62,
  input         io_iormac_63,
  input         io_iormac_64,
  input         io_iormac_65,
  input         io_iormac_66,
  input         io_iormac_67,
  input         io_iormac_68,
  input         io_iormac_69,
  input         io_iormac_70,
  input         io_iormac_71,
  input         io_iormac_72,
  input         io_iormac_73,
  input         io_iormac_74,
  input         io_iormac_75,
  input         io_iormac_76,
  input         io_iormac_77,
  input         io_iormac_78,
  input         io_iormac_79,
  input         io_iormac_80,
  input         io_iormac_81,
  input         io_iormac_82,
  input         io_iormac_83,
  input         io_iormac_84,
  input         io_iormac_85,
  input         io_iormac_86,
  input         io_iormac_87,
  input         io_iormac_88,
  input         io_iormac_89,
  input         io_iormac_90,
  input         io_iormac_91,
  input         io_iormac_92,
  input         io_iormac_93,
  input         io_iormac_94,
  input         io_iormac_95,
  input         io_iormac_96,
  input         io_iormac_97,
  input         io_iormac_98,
  input         io_iormac_99,
  input         io_iormac_100,
  input         io_iormac_101,
  input         io_iormac_102,
  input         io_iormac_103,
  input         io_iormac_104,
  input         io_iormac_105,
  input         io_iormac_106,
  input         io_iormac_107,
  input         io_iormac_108,
  input         io_iormac_109,
  input         io_iormac_110,
  input         io_iormac_111,
  input         io_iormac_112,
  input         io_iormac_113,
  input         io_iormac_114,
  input         io_iormac_115,
  input         io_iormac_116,
  input         io_iormac_117,
  input         io_iormac_118,
  input         io_iormac_119,
  input         io_iormac_120,
  input         io_iormac_121,
  input         io_iormac_122,
  input         io_iormac_123,
  input         io_iormac_124,
  input         io_iormac_125,
  input         io_iormac_126,
  input         io_iormac_127,
  input         io_iormac_128,
  input         io_iormac_129,
  input         io_iormac_130,
  input         io_iormac_131,
  input         io_iormac_132,
  input         io_iormac_133,
  input         io_iormac_134,
  input         io_iormac_135,
  input         io_iormac_136,
  input         io_iormac_137,
  input         io_iormac_138,
  input         io_iormac_139,
  input         io_iormac_140,
  input         io_iormac_141,
  input         io_iormac_142,
  input         io_iormac_143,
  input         io_iormac_144,
  input         io_iormac_145,
  input         io_iormac_146,
  input         io_iormac_147,
  input         io_iormac_148,
  input         io_iormac_149,
  input         io_iormac_150,
  input         io_iormac_151,
  input         io_iormac_152,
  input         io_iormac_153,
  input         io_iormac_154,
  input         io_iormac_155,
  input         io_iormac_156,
  input         io_iormac_157,
  input         io_iormac_158,
  input         io_iormac_159,
  input         io_iormac_160,
  input         io_iormac_161,
  input         io_iormac_162,
  input         io_iormac_163,
  input         io_iormac_164,
  input         io_iormac_165,
  input         io_iormac_166,
  input         io_iormac_167,
  input         io_iormac_168,
  input         io_iormac_169,
  input         io_iormac_170,
  input         io_iormac_171,
  input         io_iormac_172,
  input         io_iormac_173,
  input         io_iormac_174,
  input         io_iormac_175,
  input         io_iormac_176,
  input         io_iormac_177,
  input         io_iormac_178,
  input         io_iormac_179,
  input         io_iormac_180,
  input         io_iormac_181,
  input         io_iormac_182,
  input         io_iormac_183,
  input         io_iormac_184,
  input         io_iormac_185,
  input         io_iormac_186,
  input         io_iormac_187,
  input         io_iormac_188,
  input         io_iormac_189,
  input         io_iormac_190,
  input         io_iormac_191,
  input         io_iormac_192,
  input         io_iormac_193,
  input         io_iormac_194,
  input         io_iormac_195,
  input         io_iormac_196,
  input         io_iormac_197,
  input         io_iormac_198,
  input         io_iormac_199,
  input         io_iormac_200,
  input         io_iormac_201,
  input         io_iormac_202,
  input         io_iormac_203,
  input         io_iormac_204,
  input         io_iormac_205,
  input         io_iormac_206,
  input         io_iormac_207,
  input         io_iormac_208,
  input         io_iormac_209,
  input         io_iormac_210,
  input         io_iormac_211,
  input         io_iormac_212,
  input         io_iormac_213,
  input         io_iormac_214,
  input         io_iormac_215,
  input         io_iormac_216,
  input         io_iormac_217,
  input         io_iormac_218,
  input         io_iormac_219,
  input         io_iormac_220,
  input         io_iormac_221,
  input         io_iormac_222,
  input         io_iormac_223,
  input         io_iormac_224,
  input         io_iormac_225,
  input         io_iormac_226,
  input         io_iormac_227,
  input         io_iormac_228,
  input         io_iormac_229,
  input         io_iormac_230,
  input         io_iormac_231,
  input         io_iormac_232,
  input         io_iormac_233,
  input         io_iormac_234,
  input         io_iormac_235,
  input         io_iormac_236,
  input         io_iormac_237,
  input         io_iormac_238,
  input         io_iormac_239,
  input         io_iormac_240,
  input         io_iormac_241,
  input         io_iormac_242,
  input         io_iormac_243,
  input         io_iormac_244,
  input         io_iormac_245,
  input         io_iormac_246,
  input         io_iormac_247,
  input         io_iormac_248,
  input         io_iormac_249,
  input         io_iormac_250,
  input         io_iormac_251,
  input         io_iormac_252,
  input         io_iormac_253,
  input         io_iormac_254,
  input         io_iormac_255,
  output [31:0] io_out_0,
  output [31:0] io_out_1,
  output [31:0] io_out_2,
  output [31:0] io_out_3,
  output [31:0] io_out_4,
  output [31:0] io_out_5,
  output [31:0] io_out_6,
  output [31:0] io_out_7,
  output [31:0] io_out_8,
  output [31:0] io_out_9,
  output [31:0] io_out_10,
  output [31:0] io_out_11,
  output [31:0] io_out_12,
  output [31:0] io_out_13,
  output [31:0] io_out_14,
  output [31:0] io_out_15,
  output [31:0] io_out_16,
  output [31:0] io_out_17,
  output [31:0] io_out_18,
  output [31:0] io_out_19,
  output [31:0] io_out_20,
  output [31:0] io_out_21,
  output [31:0] io_out_22,
  output [31:0] io_out_23,
  output [31:0] io_out_24,
  output [31:0] io_out_25,
  output [31:0] io_out_26,
  output [31:0] io_out_27,
  output [31:0] io_out_28,
  output [31:0] io_out_29,
  output [31:0] io_out_30,
  output [31:0] io_out_31,
  output [31:0] io_out_32,
  output [31:0] io_out_33,
  output [31:0] io_out_34,
  output [31:0] io_out_35,
  output [31:0] io_out_36,
  output [31:0] io_out_37,
  output [31:0] io_out_38,
  output [31:0] io_out_39,
  output [31:0] io_out_40,
  output [31:0] io_out_41,
  output [31:0] io_out_42,
  output [31:0] io_out_43,
  output [31:0] io_out_44,
  output [31:0] io_out_45,
  output [31:0] io_out_46,
  output [31:0] io_out_47,
  output [31:0] io_out_48,
  output [31:0] io_out_49,
  output [31:0] io_out_50,
  output [31:0] io_out_51,
  output [31:0] io_out_52,
  output [31:0] io_out_53,
  output [31:0] io_out_54,
  output [31:0] io_out_55,
  output [31:0] io_out_56,
  output [31:0] io_out_57,
  output [31:0] io_out_58,
  output [31:0] io_out_59,
  output [31:0] io_out_60,
  output [31:0] io_out_61,
  output [31:0] io_out_62,
  output [31:0] io_out_63,
  output [31:0] io_out_64,
  output [31:0] io_out_65,
  output [31:0] io_out_66,
  output [31:0] io_out_67,
  output [31:0] io_out_68,
  output [31:0] io_out_69,
  output [31:0] io_out_70,
  output [31:0] io_out_71,
  output [31:0] io_out_72,
  output [31:0] io_out_73,
  output [31:0] io_out_74,
  output [31:0] io_out_75,
  output [31:0] io_out_76,
  output [31:0] io_out_77,
  output [31:0] io_out_78,
  output [31:0] io_out_79,
  output [31:0] io_out_80,
  output [31:0] io_out_81,
  output [31:0] io_out_82,
  output [31:0] io_out_83,
  output [31:0] io_out_84,
  output [31:0] io_out_85,
  output [31:0] io_out_86,
  output [31:0] io_out_87,
  output [31:0] io_out_88,
  output [31:0] io_out_89,
  output [31:0] io_out_90,
  output [31:0] io_out_91,
  output [31:0] io_out_92,
  output [31:0] io_out_93,
  output [31:0] io_out_94,
  output [31:0] io_out_95,
  output [31:0] io_out_96,
  output [31:0] io_out_97,
  output [31:0] io_out_98,
  output [31:0] io_out_99,
  output [31:0] io_out_100,
  output [31:0] io_out_101,
  output [31:0] io_out_102,
  output [31:0] io_out_103,
  output [31:0] io_out_104,
  output [31:0] io_out_105,
  output [31:0] io_out_106,
  output [31:0] io_out_107,
  output [31:0] io_out_108,
  output [31:0] io_out_109,
  output [31:0] io_out_110,
  output [31:0] io_out_111,
  output [31:0] io_out_112,
  output [31:0] io_out_113,
  output [31:0] io_out_114,
  output [31:0] io_out_115,
  output [31:0] io_out_116,
  output [31:0] io_out_117,
  output [31:0] io_out_118,
  output [31:0] io_out_119,
  output [31:0] io_out_120,
  output [31:0] io_out_121,
  output [31:0] io_out_122,
  output [31:0] io_out_123,
  output [31:0] io_out_124,
  output [31:0] io_out_125,
  output [31:0] io_out_126,
  output [31:0] io_out_127,
  output [31:0] io_out_128,
  output [31:0] io_out_129,
  output [31:0] io_out_130,
  output [31:0] io_out_131,
  output [31:0] io_out_132,
  output [31:0] io_out_133,
  output [31:0] io_out_134,
  output [31:0] io_out_135,
  output [31:0] io_out_136,
  output [31:0] io_out_137,
  output [31:0] io_out_138,
  output [31:0] io_out_139,
  output [31:0] io_out_140,
  output [31:0] io_out_141,
  output [31:0] io_out_142,
  output [31:0] io_out_143,
  output [31:0] io_out_144,
  output [31:0] io_out_145,
  output [31:0] io_out_146,
  output [31:0] io_out_147,
  output [31:0] io_out_148,
  output [31:0] io_out_149,
  output [31:0] io_out_150,
  output [31:0] io_out_151,
  output [31:0] io_out_152,
  output [31:0] io_out_153,
  output [31:0] io_out_154,
  output [31:0] io_out_155,
  output [31:0] io_out_156,
  output [31:0] io_out_157,
  output [31:0] io_out_158,
  output [31:0] io_out_159,
  output [31:0] io_out_160,
  output [31:0] io_out_161,
  output [31:0] io_out_162,
  output [31:0] io_out_163,
  output [31:0] io_out_164,
  output [31:0] io_out_165,
  output [31:0] io_out_166,
  output [31:0] io_out_167,
  output [31:0] io_out_168,
  output [31:0] io_out_169,
  output [31:0] io_out_170,
  output [31:0] io_out_171,
  output [31:0] io_out_172,
  output [31:0] io_out_173,
  output [31:0] io_out_174,
  output [31:0] io_out_175,
  output [31:0] io_out_176,
  output [31:0] io_out_177,
  output [31:0] io_out_178,
  output [31:0] io_out_179,
  output [31:0] io_out_180,
  output [31:0] io_out_181,
  output [31:0] io_out_182,
  output [31:0] io_out_183,
  output [31:0] io_out_184,
  output [31:0] io_out_185,
  output [31:0] io_out_186,
  output [31:0] io_out_187,
  output [31:0] io_out_188,
  output [31:0] io_out_189,
  output [31:0] io_out_190,
  output [31:0] io_out_191,
  output [31:0] io_out_192,
  output [31:0] io_out_193,
  output [31:0] io_out_194,
  output [31:0] io_out_195,
  output [31:0] io_out_196,
  output [31:0] io_out_197,
  output [31:0] io_out_198,
  output [31:0] io_out_199,
  output [31:0] io_out_200,
  output [31:0] io_out_201,
  output [31:0] io_out_202,
  output [31:0] io_out_203,
  output [31:0] io_out_204,
  output [31:0] io_out_205,
  output [31:0] io_out_206,
  output [31:0] io_out_207,
  output [31:0] io_out_208,
  output [31:0] io_out_209,
  output [31:0] io_out_210,
  output [31:0] io_out_211,
  output [31:0] io_out_212,
  output [31:0] io_out_213,
  output [31:0] io_out_214,
  output [31:0] io_out_215,
  output [31:0] io_out_216,
  output [31:0] io_out_217,
  output [31:0] io_out_218,
  output [31:0] io_out_219,
  output [31:0] io_out_220,
  output [31:0] io_out_221,
  output [31:0] io_out_222,
  output [31:0] io_out_223,
  output [31:0] io_out_224,
  output [31:0] io_out_225,
  output [31:0] io_out_226,
  output [31:0] io_out_227,
  output [31:0] io_out_228,
  output [31:0] io_out_229,
  output [31:0] io_out_230,
  output [31:0] io_out_231,
  output [31:0] io_out_232,
  output [31:0] io_out_233,
  output [31:0] io_out_234,
  output [31:0] io_out_235,
  output [31:0] io_out_236,
  output [31:0] io_out_237,
  output [31:0] io_out_238,
  output [31:0] io_out_239,
  output [31:0] io_out_240,
  output [31:0] io_out_241,
  output [31:0] io_out_242,
  output [31:0] io_out_243,
  output [31:0] io_out_244,
  output [31:0] io_out_245,
  output [31:0] io_out_246,
  output [31:0] io_out_247,
  output [31:0] io_out_248,
  output [31:0] io_out_249,
  output [31:0] io_out_250,
  output [31:0] io_out_251,
  output [31:0] io_out_252,
  output [31:0] io_out_253,
  output [31:0] io_out_254,
  output [31:0] io_out_255
);
  wire  bc_pe_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_1_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_1_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_1_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_2_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_2_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_2_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_2_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_2_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_2_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_2_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_2_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_2_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_3_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_3_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_3_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_3_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_3_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_3_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_3_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_3_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_3_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_4_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_4_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_4_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_4_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_4_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_4_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_4_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_4_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_4_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_5_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_5_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_5_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_5_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_5_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_5_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_5_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_5_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_5_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_6_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_6_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_6_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_6_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_6_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_6_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_6_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_6_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_6_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_7_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_7_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_7_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_7_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_7_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_7_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_7_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_7_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_7_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_8_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_8_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_8_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_8_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_8_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_8_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_8_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_8_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_8_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_9_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_9_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_9_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_9_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_9_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_9_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_9_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_9_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_9_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_10_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_10_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_10_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_10_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_10_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_10_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_10_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_10_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_10_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_11_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_11_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_11_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_11_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_11_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_11_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_11_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_11_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_11_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_12_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_12_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_12_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_12_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_12_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_12_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_12_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_12_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_12_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_13_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_13_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_13_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_13_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_13_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_13_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_13_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_13_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_13_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_14_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_14_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_14_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_14_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_14_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_14_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_14_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_14_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_14_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_15_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_15_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_15_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_15_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_15_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_15_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_15_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_15_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_15_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_16_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_16_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_16_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_16_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_16_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_16_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_16_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_16_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_16_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_17_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_17_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_17_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_17_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_17_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_17_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_17_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_17_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_17_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_18_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_18_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_18_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_18_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_18_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_18_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_18_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_18_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_18_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_19_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_19_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_19_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_19_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_19_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_19_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_19_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_19_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_19_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_20_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_20_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_20_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_20_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_20_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_20_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_20_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_20_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_20_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_21_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_21_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_21_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_21_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_21_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_21_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_21_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_21_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_21_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_22_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_22_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_22_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_22_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_22_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_22_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_22_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_22_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_22_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_23_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_23_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_23_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_23_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_23_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_23_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_23_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_23_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_23_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_24_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_24_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_24_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_24_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_24_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_24_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_24_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_24_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_24_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_25_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_25_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_25_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_25_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_25_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_25_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_25_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_25_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_25_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_26_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_26_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_26_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_26_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_26_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_26_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_26_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_26_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_26_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_27_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_27_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_27_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_27_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_27_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_27_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_27_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_27_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_27_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_28_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_28_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_28_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_28_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_28_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_28_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_28_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_28_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_28_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_29_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_29_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_29_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_29_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_29_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_29_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_29_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_29_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_29_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_30_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_30_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_30_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_30_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_30_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_30_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_30_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_30_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_30_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_31_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_31_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_31_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_31_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_31_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_31_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_31_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_31_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_31_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_32_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_32_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_32_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_32_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_32_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_32_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_32_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_32_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_32_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_33_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_33_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_33_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_33_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_33_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_33_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_33_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_33_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_33_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_34_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_34_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_34_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_34_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_34_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_34_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_34_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_34_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_34_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_35_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_35_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_35_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_35_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_35_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_35_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_35_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_35_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_35_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_36_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_36_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_36_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_36_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_36_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_36_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_36_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_36_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_36_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_37_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_37_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_37_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_37_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_37_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_37_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_37_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_37_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_37_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_38_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_38_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_38_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_38_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_38_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_38_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_38_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_38_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_38_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_39_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_39_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_39_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_39_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_39_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_39_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_39_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_39_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_39_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_40_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_40_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_40_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_40_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_40_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_40_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_40_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_40_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_40_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_41_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_41_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_41_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_41_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_41_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_41_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_41_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_41_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_41_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_42_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_42_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_42_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_42_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_42_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_42_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_42_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_42_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_42_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_43_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_43_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_43_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_43_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_43_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_43_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_43_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_43_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_43_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_44_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_44_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_44_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_44_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_44_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_44_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_44_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_44_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_44_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_45_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_45_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_45_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_45_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_45_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_45_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_45_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_45_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_45_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_46_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_46_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_46_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_46_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_46_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_46_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_46_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_46_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_46_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_47_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_47_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_47_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_47_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_47_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_47_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_47_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_47_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_47_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_48_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_48_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_48_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_48_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_48_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_48_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_48_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_48_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_48_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_49_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_49_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_49_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_49_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_49_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_49_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_49_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_49_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_49_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_50_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_50_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_50_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_50_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_50_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_50_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_50_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_50_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_50_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_51_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_51_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_51_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_51_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_51_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_51_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_51_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_51_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_51_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_52_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_52_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_52_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_52_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_52_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_52_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_52_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_52_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_52_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_53_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_53_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_53_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_53_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_53_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_53_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_53_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_53_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_53_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_54_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_54_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_54_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_54_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_54_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_54_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_54_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_54_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_54_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_55_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_55_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_55_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_55_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_55_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_55_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_55_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_55_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_55_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_56_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_56_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_56_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_56_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_56_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_56_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_56_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_56_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_56_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_57_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_57_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_57_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_57_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_57_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_57_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_57_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_57_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_57_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_58_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_58_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_58_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_58_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_58_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_58_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_58_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_58_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_58_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_59_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_59_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_59_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_59_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_59_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_59_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_59_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_59_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_59_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_60_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_60_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_60_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_60_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_60_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_60_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_60_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_60_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_60_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_61_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_61_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_61_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_61_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_61_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_61_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_61_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_61_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_61_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_62_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_62_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_62_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_62_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_62_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_62_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_62_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_62_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_62_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_63_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_63_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_63_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_63_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_63_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_63_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_63_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_63_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_63_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_64_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_64_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_64_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_64_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_64_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_64_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_64_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_64_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_64_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_65_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_65_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_65_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_65_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_65_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_65_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_65_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_65_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_65_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_66_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_66_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_66_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_66_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_66_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_66_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_66_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_66_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_66_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_67_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_67_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_67_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_67_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_67_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_67_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_67_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_67_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_67_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_68_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_68_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_68_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_68_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_68_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_68_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_68_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_68_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_68_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_69_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_69_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_69_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_69_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_69_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_69_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_69_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_69_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_69_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_70_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_70_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_70_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_70_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_70_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_70_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_70_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_70_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_70_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_71_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_71_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_71_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_71_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_71_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_71_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_71_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_71_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_71_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_72_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_72_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_72_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_72_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_72_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_72_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_72_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_72_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_72_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_73_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_73_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_73_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_73_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_73_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_73_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_73_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_73_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_73_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_74_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_74_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_74_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_74_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_74_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_74_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_74_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_74_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_74_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_75_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_75_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_75_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_75_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_75_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_75_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_75_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_75_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_75_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_76_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_76_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_76_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_76_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_76_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_76_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_76_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_76_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_76_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_77_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_77_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_77_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_77_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_77_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_77_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_77_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_77_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_77_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_78_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_78_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_78_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_78_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_78_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_78_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_78_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_78_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_78_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_79_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_79_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_79_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_79_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_79_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_79_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_79_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_79_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_79_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_80_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_80_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_80_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_80_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_80_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_80_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_80_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_80_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_80_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_81_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_81_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_81_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_81_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_81_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_81_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_81_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_81_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_81_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_82_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_82_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_82_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_82_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_82_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_82_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_82_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_82_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_82_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_83_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_83_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_83_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_83_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_83_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_83_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_83_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_83_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_83_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_84_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_84_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_84_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_84_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_84_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_84_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_84_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_84_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_84_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_85_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_85_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_85_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_85_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_85_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_85_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_85_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_85_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_85_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_86_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_86_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_86_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_86_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_86_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_86_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_86_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_86_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_86_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_87_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_87_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_87_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_87_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_87_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_87_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_87_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_87_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_87_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_88_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_88_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_88_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_88_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_88_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_88_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_88_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_88_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_88_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_89_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_89_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_89_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_89_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_89_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_89_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_89_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_89_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_89_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_90_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_90_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_90_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_90_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_90_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_90_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_90_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_90_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_90_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_91_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_91_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_91_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_91_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_91_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_91_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_91_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_91_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_91_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_92_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_92_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_92_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_92_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_92_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_92_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_92_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_92_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_92_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_93_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_93_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_93_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_93_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_93_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_93_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_93_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_93_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_93_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_94_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_94_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_94_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_94_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_94_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_94_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_94_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_94_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_94_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_95_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_95_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_95_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_95_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_95_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_95_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_95_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_95_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_95_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_96_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_96_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_96_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_96_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_96_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_96_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_96_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_96_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_96_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_97_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_97_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_97_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_97_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_97_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_97_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_97_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_97_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_97_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_98_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_98_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_98_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_98_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_98_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_98_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_98_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_98_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_98_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_99_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_99_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_99_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_99_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_99_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_99_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_99_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_99_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_99_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_100_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_100_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_100_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_100_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_100_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_100_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_100_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_100_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_100_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_101_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_101_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_101_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_101_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_101_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_101_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_101_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_101_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_101_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_102_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_102_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_102_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_102_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_102_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_102_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_102_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_102_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_102_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_103_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_103_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_103_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_103_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_103_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_103_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_103_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_103_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_103_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_104_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_104_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_104_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_104_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_104_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_104_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_104_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_104_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_104_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_105_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_105_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_105_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_105_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_105_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_105_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_105_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_105_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_105_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_106_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_106_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_106_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_106_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_106_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_106_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_106_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_106_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_106_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_107_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_107_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_107_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_107_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_107_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_107_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_107_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_107_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_107_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_108_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_108_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_108_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_108_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_108_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_108_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_108_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_108_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_108_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_109_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_109_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_109_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_109_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_109_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_109_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_109_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_109_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_109_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_110_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_110_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_110_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_110_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_110_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_110_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_110_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_110_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_110_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_111_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_111_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_111_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_111_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_111_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_111_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_111_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_111_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_111_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_112_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_112_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_112_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_112_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_112_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_112_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_112_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_112_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_112_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_113_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_113_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_113_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_113_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_113_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_113_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_113_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_113_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_113_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_114_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_114_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_114_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_114_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_114_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_114_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_114_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_114_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_114_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_115_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_115_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_115_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_115_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_115_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_115_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_115_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_115_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_115_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_116_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_116_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_116_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_116_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_116_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_116_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_116_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_116_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_116_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_117_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_117_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_117_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_117_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_117_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_117_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_117_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_117_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_117_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_118_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_118_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_118_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_118_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_118_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_118_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_118_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_118_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_118_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_119_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_119_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_119_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_119_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_119_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_119_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_119_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_119_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_119_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_120_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_120_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_120_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_120_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_120_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_120_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_120_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_120_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_120_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_121_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_121_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_121_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_121_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_121_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_121_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_121_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_121_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_121_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_122_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_122_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_122_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_122_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_122_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_122_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_122_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_122_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_122_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_123_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_123_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_123_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_123_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_123_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_123_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_123_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_123_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_123_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_124_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_124_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_124_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_124_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_124_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_124_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_124_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_124_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_124_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_125_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_125_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_125_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_125_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_125_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_125_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_125_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_125_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_125_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_126_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_126_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_126_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_126_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_126_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_126_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_126_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_126_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_126_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_127_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_127_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_127_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_127_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_127_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_127_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_127_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_127_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_127_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_128_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_128_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_128_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_128_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_128_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_128_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_128_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_128_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_128_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_129_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_129_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_129_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_129_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_129_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_129_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_129_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_129_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_129_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_130_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_130_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_130_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_130_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_130_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_130_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_130_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_130_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_130_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_131_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_131_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_131_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_131_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_131_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_131_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_131_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_131_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_131_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_132_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_132_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_132_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_132_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_132_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_132_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_132_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_132_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_132_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_133_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_133_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_133_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_133_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_133_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_133_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_133_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_133_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_133_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_134_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_134_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_134_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_134_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_134_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_134_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_134_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_134_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_134_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_135_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_135_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_135_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_135_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_135_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_135_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_135_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_135_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_135_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_136_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_136_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_136_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_136_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_136_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_136_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_136_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_136_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_136_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_137_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_137_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_137_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_137_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_137_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_137_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_137_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_137_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_137_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_138_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_138_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_138_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_138_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_138_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_138_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_138_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_138_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_138_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_139_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_139_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_139_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_139_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_139_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_139_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_139_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_139_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_139_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_140_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_140_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_140_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_140_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_140_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_140_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_140_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_140_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_140_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_141_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_141_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_141_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_141_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_141_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_141_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_141_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_141_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_141_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_142_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_142_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_142_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_142_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_142_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_142_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_142_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_142_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_142_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_143_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_143_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_143_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_143_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_143_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_143_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_143_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_143_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_143_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_144_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_144_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_144_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_144_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_144_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_144_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_144_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_144_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_144_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_145_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_145_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_145_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_145_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_145_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_145_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_145_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_145_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_145_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_146_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_146_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_146_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_146_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_146_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_146_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_146_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_146_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_146_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_147_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_147_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_147_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_147_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_147_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_147_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_147_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_147_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_147_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_148_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_148_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_148_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_148_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_148_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_148_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_148_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_148_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_148_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_149_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_149_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_149_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_149_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_149_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_149_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_149_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_149_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_149_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_150_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_150_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_150_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_150_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_150_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_150_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_150_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_150_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_150_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_151_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_151_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_151_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_151_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_151_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_151_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_151_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_151_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_151_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_152_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_152_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_152_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_152_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_152_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_152_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_152_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_152_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_152_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_153_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_153_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_153_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_153_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_153_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_153_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_153_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_153_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_153_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_154_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_154_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_154_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_154_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_154_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_154_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_154_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_154_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_154_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_155_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_155_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_155_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_155_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_155_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_155_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_155_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_155_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_155_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_156_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_156_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_156_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_156_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_156_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_156_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_156_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_156_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_156_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_157_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_157_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_157_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_157_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_157_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_157_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_157_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_157_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_157_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_158_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_158_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_158_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_158_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_158_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_158_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_158_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_158_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_158_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_159_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_159_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_159_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_159_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_159_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_159_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_159_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_159_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_159_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_160_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_160_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_160_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_160_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_160_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_160_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_160_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_160_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_160_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_161_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_161_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_161_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_161_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_161_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_161_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_161_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_161_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_161_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_162_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_162_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_162_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_162_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_162_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_162_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_162_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_162_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_162_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_163_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_163_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_163_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_163_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_163_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_163_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_163_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_163_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_163_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_164_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_164_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_164_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_164_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_164_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_164_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_164_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_164_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_164_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_165_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_165_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_165_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_165_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_165_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_165_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_165_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_165_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_165_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_166_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_166_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_166_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_166_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_166_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_166_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_166_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_166_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_166_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_167_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_167_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_167_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_167_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_167_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_167_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_167_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_167_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_167_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_168_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_168_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_168_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_168_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_168_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_168_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_168_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_168_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_168_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_169_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_169_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_169_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_169_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_169_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_169_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_169_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_169_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_169_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_170_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_170_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_170_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_170_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_170_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_170_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_170_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_170_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_170_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_171_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_171_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_171_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_171_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_171_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_171_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_171_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_171_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_171_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_172_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_172_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_172_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_172_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_172_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_172_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_172_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_172_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_172_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_173_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_173_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_173_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_173_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_173_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_173_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_173_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_173_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_173_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_174_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_174_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_174_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_174_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_174_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_174_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_174_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_174_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_174_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_175_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_175_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_175_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_175_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_175_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_175_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_175_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_175_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_175_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_176_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_176_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_176_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_176_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_176_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_176_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_176_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_176_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_176_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_177_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_177_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_177_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_177_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_177_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_177_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_177_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_177_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_177_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_178_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_178_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_178_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_178_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_178_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_178_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_178_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_178_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_178_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_179_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_179_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_179_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_179_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_179_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_179_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_179_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_179_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_179_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_180_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_180_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_180_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_180_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_180_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_180_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_180_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_180_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_180_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_181_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_181_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_181_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_181_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_181_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_181_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_181_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_181_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_181_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_182_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_182_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_182_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_182_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_182_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_182_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_182_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_182_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_182_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_183_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_183_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_183_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_183_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_183_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_183_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_183_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_183_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_183_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_184_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_184_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_184_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_184_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_184_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_184_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_184_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_184_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_184_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_185_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_185_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_185_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_185_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_185_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_185_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_185_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_185_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_185_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_186_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_186_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_186_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_186_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_186_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_186_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_186_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_186_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_186_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_187_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_187_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_187_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_187_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_187_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_187_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_187_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_187_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_187_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_188_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_188_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_188_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_188_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_188_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_188_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_188_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_188_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_188_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_189_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_189_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_189_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_189_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_189_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_189_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_189_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_189_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_189_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_190_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_190_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_190_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_190_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_190_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_190_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_190_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_190_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_190_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_191_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_191_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_191_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_191_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_191_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_191_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_191_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_191_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_191_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_192_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_192_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_192_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_192_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_192_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_192_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_192_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_192_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_192_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_193_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_193_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_193_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_193_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_193_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_193_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_193_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_193_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_193_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_194_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_194_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_194_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_194_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_194_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_194_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_194_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_194_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_194_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_195_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_195_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_195_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_195_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_195_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_195_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_195_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_195_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_195_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_196_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_196_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_196_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_196_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_196_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_196_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_196_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_196_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_196_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_197_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_197_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_197_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_197_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_197_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_197_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_197_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_197_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_197_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_198_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_198_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_198_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_198_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_198_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_198_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_198_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_198_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_198_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_199_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_199_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_199_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_199_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_199_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_199_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_199_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_199_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_199_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_200_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_200_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_200_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_200_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_200_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_200_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_200_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_200_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_200_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_201_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_201_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_201_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_201_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_201_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_201_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_201_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_201_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_201_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_202_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_202_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_202_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_202_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_202_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_202_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_202_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_202_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_202_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_203_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_203_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_203_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_203_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_203_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_203_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_203_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_203_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_203_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_204_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_204_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_204_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_204_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_204_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_204_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_204_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_204_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_204_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_205_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_205_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_205_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_205_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_205_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_205_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_205_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_205_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_205_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_206_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_206_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_206_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_206_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_206_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_206_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_206_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_206_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_206_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_207_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_207_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_207_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_207_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_207_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_207_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_207_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_207_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_207_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_208_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_208_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_208_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_208_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_208_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_208_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_208_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_208_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_208_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_209_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_209_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_209_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_209_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_209_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_209_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_209_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_209_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_209_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_210_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_210_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_210_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_210_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_210_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_210_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_210_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_210_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_210_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_211_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_211_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_211_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_211_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_211_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_211_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_211_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_211_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_211_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_212_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_212_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_212_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_212_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_212_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_212_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_212_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_212_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_212_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_213_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_213_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_213_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_213_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_213_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_213_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_213_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_213_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_213_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_214_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_214_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_214_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_214_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_214_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_214_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_214_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_214_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_214_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_215_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_215_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_215_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_215_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_215_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_215_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_215_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_215_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_215_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_216_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_216_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_216_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_216_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_216_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_216_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_216_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_216_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_216_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_217_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_217_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_217_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_217_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_217_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_217_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_217_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_217_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_217_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_218_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_218_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_218_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_218_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_218_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_218_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_218_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_218_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_218_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_219_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_219_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_219_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_219_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_219_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_219_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_219_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_219_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_219_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_220_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_220_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_220_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_220_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_220_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_220_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_220_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_220_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_220_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_221_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_221_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_221_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_221_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_221_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_221_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_221_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_221_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_221_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_222_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_222_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_222_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_222_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_222_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_222_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_222_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_222_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_222_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_223_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_223_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_223_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_223_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_223_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_223_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_223_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_223_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_223_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_224_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_224_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_224_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_224_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_224_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_224_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_224_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_224_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_224_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_225_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_225_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_225_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_225_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_225_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_225_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_225_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_225_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_225_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_226_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_226_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_226_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_226_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_226_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_226_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_226_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_226_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_226_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_227_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_227_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_227_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_227_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_227_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_227_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_227_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_227_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_227_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_228_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_228_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_228_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_228_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_228_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_228_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_228_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_228_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_228_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_229_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_229_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_229_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_229_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_229_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_229_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_229_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_229_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_229_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_230_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_230_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_230_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_230_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_230_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_230_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_230_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_230_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_230_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_231_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_231_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_231_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_231_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_231_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_231_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_231_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_231_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_231_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_232_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_232_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_232_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_232_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_232_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_232_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_232_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_232_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_232_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_233_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_233_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_233_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_233_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_233_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_233_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_233_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_233_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_233_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_234_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_234_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_234_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_234_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_234_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_234_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_234_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_234_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_234_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_235_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_235_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_235_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_235_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_235_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_235_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_235_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_235_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_235_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_236_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_236_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_236_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_236_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_236_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_236_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_236_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_236_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_236_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_237_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_237_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_237_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_237_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_237_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_237_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_237_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_237_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_237_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_238_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_238_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_238_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_238_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_238_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_238_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_238_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_238_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_238_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_239_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_239_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_239_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_239_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_239_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_239_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_239_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_239_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_239_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_240_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_240_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_240_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_240_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_240_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_240_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_240_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_240_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_240_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_241_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_241_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_241_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_241_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_241_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_241_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_241_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_241_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_241_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_242_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_242_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_242_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_242_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_242_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_242_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_242_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_242_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_242_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_243_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_243_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_243_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_243_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_243_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_243_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_243_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_243_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_243_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_244_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_244_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_244_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_244_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_244_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_244_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_244_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_244_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_244_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_245_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_245_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_245_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_245_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_245_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_245_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_245_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_245_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_245_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_246_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_246_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_246_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_246_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_246_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_246_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_246_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_246_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_246_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_247_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_247_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_247_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_247_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_247_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_247_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_247_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_247_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_247_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_248_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_248_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_248_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_248_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_248_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_248_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_248_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_248_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_248_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_249_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_249_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_249_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_249_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_249_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_249_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_249_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_249_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_249_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_250_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_250_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_250_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_250_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_250_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_250_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_250_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_250_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_250_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_251_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_251_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_251_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_251_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_251_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_251_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_251_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_251_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_251_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_252_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_252_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_252_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_252_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_252_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_252_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_252_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_252_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_252_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_253_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_253_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_253_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_253_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_253_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_253_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_253_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_253_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_253_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_254_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_254_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_254_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_254_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_254_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_254_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_254_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_254_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_254_io_res_out; // @[bc_mmul.scala 23:11]
  wire  bc_pe_255_clock; // @[bc_mmul.scala 23:11]
  wire  bc_pe_255_reset; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_255_io_ho_input; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_255_io_ve_input; // @[bc_mmul.scala 23:11]
  wire  bc_pe_255_io_input_valid; // @[bc_mmul.scala 23:11]
  wire  bc_pe_255_io_iormac; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_255_io_ve_out; // @[bc_mmul.scala 23:11]
  wire [15:0] bc_pe_255_io_ho_out; // @[bc_mmul.scala 23:11]
  wire [31:0] bc_pe_255_io_res_out; // @[bc_mmul.scala 23:11]
  bc_pe bc_pe ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_clock),
    .reset(bc_pe_reset),
    .io_ho_input(bc_pe_io_ho_input),
    .io_ve_input(bc_pe_io_ve_input),
    .io_input_valid(bc_pe_io_input_valid),
    .io_iormac(bc_pe_io_iormac),
    .io_ve_out(bc_pe_io_ve_out),
    .io_ho_out(bc_pe_io_ho_out),
    .io_res_out(bc_pe_io_res_out)
  );
  bc_pe bc_pe_1 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_1_clock),
    .reset(bc_pe_1_reset),
    .io_ho_input(bc_pe_1_io_ho_input),
    .io_ve_input(bc_pe_1_io_ve_input),
    .io_input_valid(bc_pe_1_io_input_valid),
    .io_iormac(bc_pe_1_io_iormac),
    .io_ve_out(bc_pe_1_io_ve_out),
    .io_ho_out(bc_pe_1_io_ho_out),
    .io_res_out(bc_pe_1_io_res_out)
  );
  bc_pe bc_pe_2 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_2_clock),
    .reset(bc_pe_2_reset),
    .io_ho_input(bc_pe_2_io_ho_input),
    .io_ve_input(bc_pe_2_io_ve_input),
    .io_input_valid(bc_pe_2_io_input_valid),
    .io_iormac(bc_pe_2_io_iormac),
    .io_ve_out(bc_pe_2_io_ve_out),
    .io_ho_out(bc_pe_2_io_ho_out),
    .io_res_out(bc_pe_2_io_res_out)
  );
  bc_pe bc_pe_3 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_3_clock),
    .reset(bc_pe_3_reset),
    .io_ho_input(bc_pe_3_io_ho_input),
    .io_ve_input(bc_pe_3_io_ve_input),
    .io_input_valid(bc_pe_3_io_input_valid),
    .io_iormac(bc_pe_3_io_iormac),
    .io_ve_out(bc_pe_3_io_ve_out),
    .io_ho_out(bc_pe_3_io_ho_out),
    .io_res_out(bc_pe_3_io_res_out)
  );
  bc_pe bc_pe_4 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_4_clock),
    .reset(bc_pe_4_reset),
    .io_ho_input(bc_pe_4_io_ho_input),
    .io_ve_input(bc_pe_4_io_ve_input),
    .io_input_valid(bc_pe_4_io_input_valid),
    .io_iormac(bc_pe_4_io_iormac),
    .io_ve_out(bc_pe_4_io_ve_out),
    .io_ho_out(bc_pe_4_io_ho_out),
    .io_res_out(bc_pe_4_io_res_out)
  );
  bc_pe bc_pe_5 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_5_clock),
    .reset(bc_pe_5_reset),
    .io_ho_input(bc_pe_5_io_ho_input),
    .io_ve_input(bc_pe_5_io_ve_input),
    .io_input_valid(bc_pe_5_io_input_valid),
    .io_iormac(bc_pe_5_io_iormac),
    .io_ve_out(bc_pe_5_io_ve_out),
    .io_ho_out(bc_pe_5_io_ho_out),
    .io_res_out(bc_pe_5_io_res_out)
  );
  bc_pe bc_pe_6 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_6_clock),
    .reset(bc_pe_6_reset),
    .io_ho_input(bc_pe_6_io_ho_input),
    .io_ve_input(bc_pe_6_io_ve_input),
    .io_input_valid(bc_pe_6_io_input_valid),
    .io_iormac(bc_pe_6_io_iormac),
    .io_ve_out(bc_pe_6_io_ve_out),
    .io_ho_out(bc_pe_6_io_ho_out),
    .io_res_out(bc_pe_6_io_res_out)
  );
  bc_pe bc_pe_7 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_7_clock),
    .reset(bc_pe_7_reset),
    .io_ho_input(bc_pe_7_io_ho_input),
    .io_ve_input(bc_pe_7_io_ve_input),
    .io_input_valid(bc_pe_7_io_input_valid),
    .io_iormac(bc_pe_7_io_iormac),
    .io_ve_out(bc_pe_7_io_ve_out),
    .io_ho_out(bc_pe_7_io_ho_out),
    .io_res_out(bc_pe_7_io_res_out)
  );
  bc_pe bc_pe_8 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_8_clock),
    .reset(bc_pe_8_reset),
    .io_ho_input(bc_pe_8_io_ho_input),
    .io_ve_input(bc_pe_8_io_ve_input),
    .io_input_valid(bc_pe_8_io_input_valid),
    .io_iormac(bc_pe_8_io_iormac),
    .io_ve_out(bc_pe_8_io_ve_out),
    .io_ho_out(bc_pe_8_io_ho_out),
    .io_res_out(bc_pe_8_io_res_out)
  );
  bc_pe bc_pe_9 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_9_clock),
    .reset(bc_pe_9_reset),
    .io_ho_input(bc_pe_9_io_ho_input),
    .io_ve_input(bc_pe_9_io_ve_input),
    .io_input_valid(bc_pe_9_io_input_valid),
    .io_iormac(bc_pe_9_io_iormac),
    .io_ve_out(bc_pe_9_io_ve_out),
    .io_ho_out(bc_pe_9_io_ho_out),
    .io_res_out(bc_pe_9_io_res_out)
  );
  bc_pe bc_pe_10 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_10_clock),
    .reset(bc_pe_10_reset),
    .io_ho_input(bc_pe_10_io_ho_input),
    .io_ve_input(bc_pe_10_io_ve_input),
    .io_input_valid(bc_pe_10_io_input_valid),
    .io_iormac(bc_pe_10_io_iormac),
    .io_ve_out(bc_pe_10_io_ve_out),
    .io_ho_out(bc_pe_10_io_ho_out),
    .io_res_out(bc_pe_10_io_res_out)
  );
  bc_pe bc_pe_11 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_11_clock),
    .reset(bc_pe_11_reset),
    .io_ho_input(bc_pe_11_io_ho_input),
    .io_ve_input(bc_pe_11_io_ve_input),
    .io_input_valid(bc_pe_11_io_input_valid),
    .io_iormac(bc_pe_11_io_iormac),
    .io_ve_out(bc_pe_11_io_ve_out),
    .io_ho_out(bc_pe_11_io_ho_out),
    .io_res_out(bc_pe_11_io_res_out)
  );
  bc_pe bc_pe_12 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_12_clock),
    .reset(bc_pe_12_reset),
    .io_ho_input(bc_pe_12_io_ho_input),
    .io_ve_input(bc_pe_12_io_ve_input),
    .io_input_valid(bc_pe_12_io_input_valid),
    .io_iormac(bc_pe_12_io_iormac),
    .io_ve_out(bc_pe_12_io_ve_out),
    .io_ho_out(bc_pe_12_io_ho_out),
    .io_res_out(bc_pe_12_io_res_out)
  );
  bc_pe bc_pe_13 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_13_clock),
    .reset(bc_pe_13_reset),
    .io_ho_input(bc_pe_13_io_ho_input),
    .io_ve_input(bc_pe_13_io_ve_input),
    .io_input_valid(bc_pe_13_io_input_valid),
    .io_iormac(bc_pe_13_io_iormac),
    .io_ve_out(bc_pe_13_io_ve_out),
    .io_ho_out(bc_pe_13_io_ho_out),
    .io_res_out(bc_pe_13_io_res_out)
  );
  bc_pe bc_pe_14 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_14_clock),
    .reset(bc_pe_14_reset),
    .io_ho_input(bc_pe_14_io_ho_input),
    .io_ve_input(bc_pe_14_io_ve_input),
    .io_input_valid(bc_pe_14_io_input_valid),
    .io_iormac(bc_pe_14_io_iormac),
    .io_ve_out(bc_pe_14_io_ve_out),
    .io_ho_out(bc_pe_14_io_ho_out),
    .io_res_out(bc_pe_14_io_res_out)
  );
  bc_pe bc_pe_15 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_15_clock),
    .reset(bc_pe_15_reset),
    .io_ho_input(bc_pe_15_io_ho_input),
    .io_ve_input(bc_pe_15_io_ve_input),
    .io_input_valid(bc_pe_15_io_input_valid),
    .io_iormac(bc_pe_15_io_iormac),
    .io_ve_out(bc_pe_15_io_ve_out),
    .io_ho_out(bc_pe_15_io_ho_out),
    .io_res_out(bc_pe_15_io_res_out)
  );
  bc_pe bc_pe_16 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_16_clock),
    .reset(bc_pe_16_reset),
    .io_ho_input(bc_pe_16_io_ho_input),
    .io_ve_input(bc_pe_16_io_ve_input),
    .io_input_valid(bc_pe_16_io_input_valid),
    .io_iormac(bc_pe_16_io_iormac),
    .io_ve_out(bc_pe_16_io_ve_out),
    .io_ho_out(bc_pe_16_io_ho_out),
    .io_res_out(bc_pe_16_io_res_out)
  );
  bc_pe bc_pe_17 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_17_clock),
    .reset(bc_pe_17_reset),
    .io_ho_input(bc_pe_17_io_ho_input),
    .io_ve_input(bc_pe_17_io_ve_input),
    .io_input_valid(bc_pe_17_io_input_valid),
    .io_iormac(bc_pe_17_io_iormac),
    .io_ve_out(bc_pe_17_io_ve_out),
    .io_ho_out(bc_pe_17_io_ho_out),
    .io_res_out(bc_pe_17_io_res_out)
  );
  bc_pe bc_pe_18 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_18_clock),
    .reset(bc_pe_18_reset),
    .io_ho_input(bc_pe_18_io_ho_input),
    .io_ve_input(bc_pe_18_io_ve_input),
    .io_input_valid(bc_pe_18_io_input_valid),
    .io_iormac(bc_pe_18_io_iormac),
    .io_ve_out(bc_pe_18_io_ve_out),
    .io_ho_out(bc_pe_18_io_ho_out),
    .io_res_out(bc_pe_18_io_res_out)
  );
  bc_pe bc_pe_19 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_19_clock),
    .reset(bc_pe_19_reset),
    .io_ho_input(bc_pe_19_io_ho_input),
    .io_ve_input(bc_pe_19_io_ve_input),
    .io_input_valid(bc_pe_19_io_input_valid),
    .io_iormac(bc_pe_19_io_iormac),
    .io_ve_out(bc_pe_19_io_ve_out),
    .io_ho_out(bc_pe_19_io_ho_out),
    .io_res_out(bc_pe_19_io_res_out)
  );
  bc_pe bc_pe_20 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_20_clock),
    .reset(bc_pe_20_reset),
    .io_ho_input(bc_pe_20_io_ho_input),
    .io_ve_input(bc_pe_20_io_ve_input),
    .io_input_valid(bc_pe_20_io_input_valid),
    .io_iormac(bc_pe_20_io_iormac),
    .io_ve_out(bc_pe_20_io_ve_out),
    .io_ho_out(bc_pe_20_io_ho_out),
    .io_res_out(bc_pe_20_io_res_out)
  );
  bc_pe bc_pe_21 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_21_clock),
    .reset(bc_pe_21_reset),
    .io_ho_input(bc_pe_21_io_ho_input),
    .io_ve_input(bc_pe_21_io_ve_input),
    .io_input_valid(bc_pe_21_io_input_valid),
    .io_iormac(bc_pe_21_io_iormac),
    .io_ve_out(bc_pe_21_io_ve_out),
    .io_ho_out(bc_pe_21_io_ho_out),
    .io_res_out(bc_pe_21_io_res_out)
  );
  bc_pe bc_pe_22 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_22_clock),
    .reset(bc_pe_22_reset),
    .io_ho_input(bc_pe_22_io_ho_input),
    .io_ve_input(bc_pe_22_io_ve_input),
    .io_input_valid(bc_pe_22_io_input_valid),
    .io_iormac(bc_pe_22_io_iormac),
    .io_ve_out(bc_pe_22_io_ve_out),
    .io_ho_out(bc_pe_22_io_ho_out),
    .io_res_out(bc_pe_22_io_res_out)
  );
  bc_pe bc_pe_23 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_23_clock),
    .reset(bc_pe_23_reset),
    .io_ho_input(bc_pe_23_io_ho_input),
    .io_ve_input(bc_pe_23_io_ve_input),
    .io_input_valid(bc_pe_23_io_input_valid),
    .io_iormac(bc_pe_23_io_iormac),
    .io_ve_out(bc_pe_23_io_ve_out),
    .io_ho_out(bc_pe_23_io_ho_out),
    .io_res_out(bc_pe_23_io_res_out)
  );
  bc_pe bc_pe_24 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_24_clock),
    .reset(bc_pe_24_reset),
    .io_ho_input(bc_pe_24_io_ho_input),
    .io_ve_input(bc_pe_24_io_ve_input),
    .io_input_valid(bc_pe_24_io_input_valid),
    .io_iormac(bc_pe_24_io_iormac),
    .io_ve_out(bc_pe_24_io_ve_out),
    .io_ho_out(bc_pe_24_io_ho_out),
    .io_res_out(bc_pe_24_io_res_out)
  );
  bc_pe bc_pe_25 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_25_clock),
    .reset(bc_pe_25_reset),
    .io_ho_input(bc_pe_25_io_ho_input),
    .io_ve_input(bc_pe_25_io_ve_input),
    .io_input_valid(bc_pe_25_io_input_valid),
    .io_iormac(bc_pe_25_io_iormac),
    .io_ve_out(bc_pe_25_io_ve_out),
    .io_ho_out(bc_pe_25_io_ho_out),
    .io_res_out(bc_pe_25_io_res_out)
  );
  bc_pe bc_pe_26 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_26_clock),
    .reset(bc_pe_26_reset),
    .io_ho_input(bc_pe_26_io_ho_input),
    .io_ve_input(bc_pe_26_io_ve_input),
    .io_input_valid(bc_pe_26_io_input_valid),
    .io_iormac(bc_pe_26_io_iormac),
    .io_ve_out(bc_pe_26_io_ve_out),
    .io_ho_out(bc_pe_26_io_ho_out),
    .io_res_out(bc_pe_26_io_res_out)
  );
  bc_pe bc_pe_27 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_27_clock),
    .reset(bc_pe_27_reset),
    .io_ho_input(bc_pe_27_io_ho_input),
    .io_ve_input(bc_pe_27_io_ve_input),
    .io_input_valid(bc_pe_27_io_input_valid),
    .io_iormac(bc_pe_27_io_iormac),
    .io_ve_out(bc_pe_27_io_ve_out),
    .io_ho_out(bc_pe_27_io_ho_out),
    .io_res_out(bc_pe_27_io_res_out)
  );
  bc_pe bc_pe_28 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_28_clock),
    .reset(bc_pe_28_reset),
    .io_ho_input(bc_pe_28_io_ho_input),
    .io_ve_input(bc_pe_28_io_ve_input),
    .io_input_valid(bc_pe_28_io_input_valid),
    .io_iormac(bc_pe_28_io_iormac),
    .io_ve_out(bc_pe_28_io_ve_out),
    .io_ho_out(bc_pe_28_io_ho_out),
    .io_res_out(bc_pe_28_io_res_out)
  );
  bc_pe bc_pe_29 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_29_clock),
    .reset(bc_pe_29_reset),
    .io_ho_input(bc_pe_29_io_ho_input),
    .io_ve_input(bc_pe_29_io_ve_input),
    .io_input_valid(bc_pe_29_io_input_valid),
    .io_iormac(bc_pe_29_io_iormac),
    .io_ve_out(bc_pe_29_io_ve_out),
    .io_ho_out(bc_pe_29_io_ho_out),
    .io_res_out(bc_pe_29_io_res_out)
  );
  bc_pe bc_pe_30 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_30_clock),
    .reset(bc_pe_30_reset),
    .io_ho_input(bc_pe_30_io_ho_input),
    .io_ve_input(bc_pe_30_io_ve_input),
    .io_input_valid(bc_pe_30_io_input_valid),
    .io_iormac(bc_pe_30_io_iormac),
    .io_ve_out(bc_pe_30_io_ve_out),
    .io_ho_out(bc_pe_30_io_ho_out),
    .io_res_out(bc_pe_30_io_res_out)
  );
  bc_pe bc_pe_31 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_31_clock),
    .reset(bc_pe_31_reset),
    .io_ho_input(bc_pe_31_io_ho_input),
    .io_ve_input(bc_pe_31_io_ve_input),
    .io_input_valid(bc_pe_31_io_input_valid),
    .io_iormac(bc_pe_31_io_iormac),
    .io_ve_out(bc_pe_31_io_ve_out),
    .io_ho_out(bc_pe_31_io_ho_out),
    .io_res_out(bc_pe_31_io_res_out)
  );
  bc_pe bc_pe_32 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_32_clock),
    .reset(bc_pe_32_reset),
    .io_ho_input(bc_pe_32_io_ho_input),
    .io_ve_input(bc_pe_32_io_ve_input),
    .io_input_valid(bc_pe_32_io_input_valid),
    .io_iormac(bc_pe_32_io_iormac),
    .io_ve_out(bc_pe_32_io_ve_out),
    .io_ho_out(bc_pe_32_io_ho_out),
    .io_res_out(bc_pe_32_io_res_out)
  );
  bc_pe bc_pe_33 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_33_clock),
    .reset(bc_pe_33_reset),
    .io_ho_input(bc_pe_33_io_ho_input),
    .io_ve_input(bc_pe_33_io_ve_input),
    .io_input_valid(bc_pe_33_io_input_valid),
    .io_iormac(bc_pe_33_io_iormac),
    .io_ve_out(bc_pe_33_io_ve_out),
    .io_ho_out(bc_pe_33_io_ho_out),
    .io_res_out(bc_pe_33_io_res_out)
  );
  bc_pe bc_pe_34 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_34_clock),
    .reset(bc_pe_34_reset),
    .io_ho_input(bc_pe_34_io_ho_input),
    .io_ve_input(bc_pe_34_io_ve_input),
    .io_input_valid(bc_pe_34_io_input_valid),
    .io_iormac(bc_pe_34_io_iormac),
    .io_ve_out(bc_pe_34_io_ve_out),
    .io_ho_out(bc_pe_34_io_ho_out),
    .io_res_out(bc_pe_34_io_res_out)
  );
  bc_pe bc_pe_35 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_35_clock),
    .reset(bc_pe_35_reset),
    .io_ho_input(bc_pe_35_io_ho_input),
    .io_ve_input(bc_pe_35_io_ve_input),
    .io_input_valid(bc_pe_35_io_input_valid),
    .io_iormac(bc_pe_35_io_iormac),
    .io_ve_out(bc_pe_35_io_ve_out),
    .io_ho_out(bc_pe_35_io_ho_out),
    .io_res_out(bc_pe_35_io_res_out)
  );
  bc_pe bc_pe_36 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_36_clock),
    .reset(bc_pe_36_reset),
    .io_ho_input(bc_pe_36_io_ho_input),
    .io_ve_input(bc_pe_36_io_ve_input),
    .io_input_valid(bc_pe_36_io_input_valid),
    .io_iormac(bc_pe_36_io_iormac),
    .io_ve_out(bc_pe_36_io_ve_out),
    .io_ho_out(bc_pe_36_io_ho_out),
    .io_res_out(bc_pe_36_io_res_out)
  );
  bc_pe bc_pe_37 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_37_clock),
    .reset(bc_pe_37_reset),
    .io_ho_input(bc_pe_37_io_ho_input),
    .io_ve_input(bc_pe_37_io_ve_input),
    .io_input_valid(bc_pe_37_io_input_valid),
    .io_iormac(bc_pe_37_io_iormac),
    .io_ve_out(bc_pe_37_io_ve_out),
    .io_ho_out(bc_pe_37_io_ho_out),
    .io_res_out(bc_pe_37_io_res_out)
  );
  bc_pe bc_pe_38 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_38_clock),
    .reset(bc_pe_38_reset),
    .io_ho_input(bc_pe_38_io_ho_input),
    .io_ve_input(bc_pe_38_io_ve_input),
    .io_input_valid(bc_pe_38_io_input_valid),
    .io_iormac(bc_pe_38_io_iormac),
    .io_ve_out(bc_pe_38_io_ve_out),
    .io_ho_out(bc_pe_38_io_ho_out),
    .io_res_out(bc_pe_38_io_res_out)
  );
  bc_pe bc_pe_39 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_39_clock),
    .reset(bc_pe_39_reset),
    .io_ho_input(bc_pe_39_io_ho_input),
    .io_ve_input(bc_pe_39_io_ve_input),
    .io_input_valid(bc_pe_39_io_input_valid),
    .io_iormac(bc_pe_39_io_iormac),
    .io_ve_out(bc_pe_39_io_ve_out),
    .io_ho_out(bc_pe_39_io_ho_out),
    .io_res_out(bc_pe_39_io_res_out)
  );
  bc_pe bc_pe_40 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_40_clock),
    .reset(bc_pe_40_reset),
    .io_ho_input(bc_pe_40_io_ho_input),
    .io_ve_input(bc_pe_40_io_ve_input),
    .io_input_valid(bc_pe_40_io_input_valid),
    .io_iormac(bc_pe_40_io_iormac),
    .io_ve_out(bc_pe_40_io_ve_out),
    .io_ho_out(bc_pe_40_io_ho_out),
    .io_res_out(bc_pe_40_io_res_out)
  );
  bc_pe bc_pe_41 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_41_clock),
    .reset(bc_pe_41_reset),
    .io_ho_input(bc_pe_41_io_ho_input),
    .io_ve_input(bc_pe_41_io_ve_input),
    .io_input_valid(bc_pe_41_io_input_valid),
    .io_iormac(bc_pe_41_io_iormac),
    .io_ve_out(bc_pe_41_io_ve_out),
    .io_ho_out(bc_pe_41_io_ho_out),
    .io_res_out(bc_pe_41_io_res_out)
  );
  bc_pe bc_pe_42 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_42_clock),
    .reset(bc_pe_42_reset),
    .io_ho_input(bc_pe_42_io_ho_input),
    .io_ve_input(bc_pe_42_io_ve_input),
    .io_input_valid(bc_pe_42_io_input_valid),
    .io_iormac(bc_pe_42_io_iormac),
    .io_ve_out(bc_pe_42_io_ve_out),
    .io_ho_out(bc_pe_42_io_ho_out),
    .io_res_out(bc_pe_42_io_res_out)
  );
  bc_pe bc_pe_43 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_43_clock),
    .reset(bc_pe_43_reset),
    .io_ho_input(bc_pe_43_io_ho_input),
    .io_ve_input(bc_pe_43_io_ve_input),
    .io_input_valid(bc_pe_43_io_input_valid),
    .io_iormac(bc_pe_43_io_iormac),
    .io_ve_out(bc_pe_43_io_ve_out),
    .io_ho_out(bc_pe_43_io_ho_out),
    .io_res_out(bc_pe_43_io_res_out)
  );
  bc_pe bc_pe_44 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_44_clock),
    .reset(bc_pe_44_reset),
    .io_ho_input(bc_pe_44_io_ho_input),
    .io_ve_input(bc_pe_44_io_ve_input),
    .io_input_valid(bc_pe_44_io_input_valid),
    .io_iormac(bc_pe_44_io_iormac),
    .io_ve_out(bc_pe_44_io_ve_out),
    .io_ho_out(bc_pe_44_io_ho_out),
    .io_res_out(bc_pe_44_io_res_out)
  );
  bc_pe bc_pe_45 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_45_clock),
    .reset(bc_pe_45_reset),
    .io_ho_input(bc_pe_45_io_ho_input),
    .io_ve_input(bc_pe_45_io_ve_input),
    .io_input_valid(bc_pe_45_io_input_valid),
    .io_iormac(bc_pe_45_io_iormac),
    .io_ve_out(bc_pe_45_io_ve_out),
    .io_ho_out(bc_pe_45_io_ho_out),
    .io_res_out(bc_pe_45_io_res_out)
  );
  bc_pe bc_pe_46 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_46_clock),
    .reset(bc_pe_46_reset),
    .io_ho_input(bc_pe_46_io_ho_input),
    .io_ve_input(bc_pe_46_io_ve_input),
    .io_input_valid(bc_pe_46_io_input_valid),
    .io_iormac(bc_pe_46_io_iormac),
    .io_ve_out(bc_pe_46_io_ve_out),
    .io_ho_out(bc_pe_46_io_ho_out),
    .io_res_out(bc_pe_46_io_res_out)
  );
  bc_pe bc_pe_47 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_47_clock),
    .reset(bc_pe_47_reset),
    .io_ho_input(bc_pe_47_io_ho_input),
    .io_ve_input(bc_pe_47_io_ve_input),
    .io_input_valid(bc_pe_47_io_input_valid),
    .io_iormac(bc_pe_47_io_iormac),
    .io_ve_out(bc_pe_47_io_ve_out),
    .io_ho_out(bc_pe_47_io_ho_out),
    .io_res_out(bc_pe_47_io_res_out)
  );
  bc_pe bc_pe_48 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_48_clock),
    .reset(bc_pe_48_reset),
    .io_ho_input(bc_pe_48_io_ho_input),
    .io_ve_input(bc_pe_48_io_ve_input),
    .io_input_valid(bc_pe_48_io_input_valid),
    .io_iormac(bc_pe_48_io_iormac),
    .io_ve_out(bc_pe_48_io_ve_out),
    .io_ho_out(bc_pe_48_io_ho_out),
    .io_res_out(bc_pe_48_io_res_out)
  );
  bc_pe bc_pe_49 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_49_clock),
    .reset(bc_pe_49_reset),
    .io_ho_input(bc_pe_49_io_ho_input),
    .io_ve_input(bc_pe_49_io_ve_input),
    .io_input_valid(bc_pe_49_io_input_valid),
    .io_iormac(bc_pe_49_io_iormac),
    .io_ve_out(bc_pe_49_io_ve_out),
    .io_ho_out(bc_pe_49_io_ho_out),
    .io_res_out(bc_pe_49_io_res_out)
  );
  bc_pe bc_pe_50 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_50_clock),
    .reset(bc_pe_50_reset),
    .io_ho_input(bc_pe_50_io_ho_input),
    .io_ve_input(bc_pe_50_io_ve_input),
    .io_input_valid(bc_pe_50_io_input_valid),
    .io_iormac(bc_pe_50_io_iormac),
    .io_ve_out(bc_pe_50_io_ve_out),
    .io_ho_out(bc_pe_50_io_ho_out),
    .io_res_out(bc_pe_50_io_res_out)
  );
  bc_pe bc_pe_51 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_51_clock),
    .reset(bc_pe_51_reset),
    .io_ho_input(bc_pe_51_io_ho_input),
    .io_ve_input(bc_pe_51_io_ve_input),
    .io_input_valid(bc_pe_51_io_input_valid),
    .io_iormac(bc_pe_51_io_iormac),
    .io_ve_out(bc_pe_51_io_ve_out),
    .io_ho_out(bc_pe_51_io_ho_out),
    .io_res_out(bc_pe_51_io_res_out)
  );
  bc_pe bc_pe_52 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_52_clock),
    .reset(bc_pe_52_reset),
    .io_ho_input(bc_pe_52_io_ho_input),
    .io_ve_input(bc_pe_52_io_ve_input),
    .io_input_valid(bc_pe_52_io_input_valid),
    .io_iormac(bc_pe_52_io_iormac),
    .io_ve_out(bc_pe_52_io_ve_out),
    .io_ho_out(bc_pe_52_io_ho_out),
    .io_res_out(bc_pe_52_io_res_out)
  );
  bc_pe bc_pe_53 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_53_clock),
    .reset(bc_pe_53_reset),
    .io_ho_input(bc_pe_53_io_ho_input),
    .io_ve_input(bc_pe_53_io_ve_input),
    .io_input_valid(bc_pe_53_io_input_valid),
    .io_iormac(bc_pe_53_io_iormac),
    .io_ve_out(bc_pe_53_io_ve_out),
    .io_ho_out(bc_pe_53_io_ho_out),
    .io_res_out(bc_pe_53_io_res_out)
  );
  bc_pe bc_pe_54 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_54_clock),
    .reset(bc_pe_54_reset),
    .io_ho_input(bc_pe_54_io_ho_input),
    .io_ve_input(bc_pe_54_io_ve_input),
    .io_input_valid(bc_pe_54_io_input_valid),
    .io_iormac(bc_pe_54_io_iormac),
    .io_ve_out(bc_pe_54_io_ve_out),
    .io_ho_out(bc_pe_54_io_ho_out),
    .io_res_out(bc_pe_54_io_res_out)
  );
  bc_pe bc_pe_55 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_55_clock),
    .reset(bc_pe_55_reset),
    .io_ho_input(bc_pe_55_io_ho_input),
    .io_ve_input(bc_pe_55_io_ve_input),
    .io_input_valid(bc_pe_55_io_input_valid),
    .io_iormac(bc_pe_55_io_iormac),
    .io_ve_out(bc_pe_55_io_ve_out),
    .io_ho_out(bc_pe_55_io_ho_out),
    .io_res_out(bc_pe_55_io_res_out)
  );
  bc_pe bc_pe_56 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_56_clock),
    .reset(bc_pe_56_reset),
    .io_ho_input(bc_pe_56_io_ho_input),
    .io_ve_input(bc_pe_56_io_ve_input),
    .io_input_valid(bc_pe_56_io_input_valid),
    .io_iormac(bc_pe_56_io_iormac),
    .io_ve_out(bc_pe_56_io_ve_out),
    .io_ho_out(bc_pe_56_io_ho_out),
    .io_res_out(bc_pe_56_io_res_out)
  );
  bc_pe bc_pe_57 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_57_clock),
    .reset(bc_pe_57_reset),
    .io_ho_input(bc_pe_57_io_ho_input),
    .io_ve_input(bc_pe_57_io_ve_input),
    .io_input_valid(bc_pe_57_io_input_valid),
    .io_iormac(bc_pe_57_io_iormac),
    .io_ve_out(bc_pe_57_io_ve_out),
    .io_ho_out(bc_pe_57_io_ho_out),
    .io_res_out(bc_pe_57_io_res_out)
  );
  bc_pe bc_pe_58 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_58_clock),
    .reset(bc_pe_58_reset),
    .io_ho_input(bc_pe_58_io_ho_input),
    .io_ve_input(bc_pe_58_io_ve_input),
    .io_input_valid(bc_pe_58_io_input_valid),
    .io_iormac(bc_pe_58_io_iormac),
    .io_ve_out(bc_pe_58_io_ve_out),
    .io_ho_out(bc_pe_58_io_ho_out),
    .io_res_out(bc_pe_58_io_res_out)
  );
  bc_pe bc_pe_59 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_59_clock),
    .reset(bc_pe_59_reset),
    .io_ho_input(bc_pe_59_io_ho_input),
    .io_ve_input(bc_pe_59_io_ve_input),
    .io_input_valid(bc_pe_59_io_input_valid),
    .io_iormac(bc_pe_59_io_iormac),
    .io_ve_out(bc_pe_59_io_ve_out),
    .io_ho_out(bc_pe_59_io_ho_out),
    .io_res_out(bc_pe_59_io_res_out)
  );
  bc_pe bc_pe_60 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_60_clock),
    .reset(bc_pe_60_reset),
    .io_ho_input(bc_pe_60_io_ho_input),
    .io_ve_input(bc_pe_60_io_ve_input),
    .io_input_valid(bc_pe_60_io_input_valid),
    .io_iormac(bc_pe_60_io_iormac),
    .io_ve_out(bc_pe_60_io_ve_out),
    .io_ho_out(bc_pe_60_io_ho_out),
    .io_res_out(bc_pe_60_io_res_out)
  );
  bc_pe bc_pe_61 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_61_clock),
    .reset(bc_pe_61_reset),
    .io_ho_input(bc_pe_61_io_ho_input),
    .io_ve_input(bc_pe_61_io_ve_input),
    .io_input_valid(bc_pe_61_io_input_valid),
    .io_iormac(bc_pe_61_io_iormac),
    .io_ve_out(bc_pe_61_io_ve_out),
    .io_ho_out(bc_pe_61_io_ho_out),
    .io_res_out(bc_pe_61_io_res_out)
  );
  bc_pe bc_pe_62 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_62_clock),
    .reset(bc_pe_62_reset),
    .io_ho_input(bc_pe_62_io_ho_input),
    .io_ve_input(bc_pe_62_io_ve_input),
    .io_input_valid(bc_pe_62_io_input_valid),
    .io_iormac(bc_pe_62_io_iormac),
    .io_ve_out(bc_pe_62_io_ve_out),
    .io_ho_out(bc_pe_62_io_ho_out),
    .io_res_out(bc_pe_62_io_res_out)
  );
  bc_pe bc_pe_63 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_63_clock),
    .reset(bc_pe_63_reset),
    .io_ho_input(bc_pe_63_io_ho_input),
    .io_ve_input(bc_pe_63_io_ve_input),
    .io_input_valid(bc_pe_63_io_input_valid),
    .io_iormac(bc_pe_63_io_iormac),
    .io_ve_out(bc_pe_63_io_ve_out),
    .io_ho_out(bc_pe_63_io_ho_out),
    .io_res_out(bc_pe_63_io_res_out)
  );
  bc_pe bc_pe_64 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_64_clock),
    .reset(bc_pe_64_reset),
    .io_ho_input(bc_pe_64_io_ho_input),
    .io_ve_input(bc_pe_64_io_ve_input),
    .io_input_valid(bc_pe_64_io_input_valid),
    .io_iormac(bc_pe_64_io_iormac),
    .io_ve_out(bc_pe_64_io_ve_out),
    .io_ho_out(bc_pe_64_io_ho_out),
    .io_res_out(bc_pe_64_io_res_out)
  );
  bc_pe bc_pe_65 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_65_clock),
    .reset(bc_pe_65_reset),
    .io_ho_input(bc_pe_65_io_ho_input),
    .io_ve_input(bc_pe_65_io_ve_input),
    .io_input_valid(bc_pe_65_io_input_valid),
    .io_iormac(bc_pe_65_io_iormac),
    .io_ve_out(bc_pe_65_io_ve_out),
    .io_ho_out(bc_pe_65_io_ho_out),
    .io_res_out(bc_pe_65_io_res_out)
  );
  bc_pe bc_pe_66 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_66_clock),
    .reset(bc_pe_66_reset),
    .io_ho_input(bc_pe_66_io_ho_input),
    .io_ve_input(bc_pe_66_io_ve_input),
    .io_input_valid(bc_pe_66_io_input_valid),
    .io_iormac(bc_pe_66_io_iormac),
    .io_ve_out(bc_pe_66_io_ve_out),
    .io_ho_out(bc_pe_66_io_ho_out),
    .io_res_out(bc_pe_66_io_res_out)
  );
  bc_pe bc_pe_67 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_67_clock),
    .reset(bc_pe_67_reset),
    .io_ho_input(bc_pe_67_io_ho_input),
    .io_ve_input(bc_pe_67_io_ve_input),
    .io_input_valid(bc_pe_67_io_input_valid),
    .io_iormac(bc_pe_67_io_iormac),
    .io_ve_out(bc_pe_67_io_ve_out),
    .io_ho_out(bc_pe_67_io_ho_out),
    .io_res_out(bc_pe_67_io_res_out)
  );
  bc_pe bc_pe_68 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_68_clock),
    .reset(bc_pe_68_reset),
    .io_ho_input(bc_pe_68_io_ho_input),
    .io_ve_input(bc_pe_68_io_ve_input),
    .io_input_valid(bc_pe_68_io_input_valid),
    .io_iormac(bc_pe_68_io_iormac),
    .io_ve_out(bc_pe_68_io_ve_out),
    .io_ho_out(bc_pe_68_io_ho_out),
    .io_res_out(bc_pe_68_io_res_out)
  );
  bc_pe bc_pe_69 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_69_clock),
    .reset(bc_pe_69_reset),
    .io_ho_input(bc_pe_69_io_ho_input),
    .io_ve_input(bc_pe_69_io_ve_input),
    .io_input_valid(bc_pe_69_io_input_valid),
    .io_iormac(bc_pe_69_io_iormac),
    .io_ve_out(bc_pe_69_io_ve_out),
    .io_ho_out(bc_pe_69_io_ho_out),
    .io_res_out(bc_pe_69_io_res_out)
  );
  bc_pe bc_pe_70 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_70_clock),
    .reset(bc_pe_70_reset),
    .io_ho_input(bc_pe_70_io_ho_input),
    .io_ve_input(bc_pe_70_io_ve_input),
    .io_input_valid(bc_pe_70_io_input_valid),
    .io_iormac(bc_pe_70_io_iormac),
    .io_ve_out(bc_pe_70_io_ve_out),
    .io_ho_out(bc_pe_70_io_ho_out),
    .io_res_out(bc_pe_70_io_res_out)
  );
  bc_pe bc_pe_71 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_71_clock),
    .reset(bc_pe_71_reset),
    .io_ho_input(bc_pe_71_io_ho_input),
    .io_ve_input(bc_pe_71_io_ve_input),
    .io_input_valid(bc_pe_71_io_input_valid),
    .io_iormac(bc_pe_71_io_iormac),
    .io_ve_out(bc_pe_71_io_ve_out),
    .io_ho_out(bc_pe_71_io_ho_out),
    .io_res_out(bc_pe_71_io_res_out)
  );
  bc_pe bc_pe_72 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_72_clock),
    .reset(bc_pe_72_reset),
    .io_ho_input(bc_pe_72_io_ho_input),
    .io_ve_input(bc_pe_72_io_ve_input),
    .io_input_valid(bc_pe_72_io_input_valid),
    .io_iormac(bc_pe_72_io_iormac),
    .io_ve_out(bc_pe_72_io_ve_out),
    .io_ho_out(bc_pe_72_io_ho_out),
    .io_res_out(bc_pe_72_io_res_out)
  );
  bc_pe bc_pe_73 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_73_clock),
    .reset(bc_pe_73_reset),
    .io_ho_input(bc_pe_73_io_ho_input),
    .io_ve_input(bc_pe_73_io_ve_input),
    .io_input_valid(bc_pe_73_io_input_valid),
    .io_iormac(bc_pe_73_io_iormac),
    .io_ve_out(bc_pe_73_io_ve_out),
    .io_ho_out(bc_pe_73_io_ho_out),
    .io_res_out(bc_pe_73_io_res_out)
  );
  bc_pe bc_pe_74 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_74_clock),
    .reset(bc_pe_74_reset),
    .io_ho_input(bc_pe_74_io_ho_input),
    .io_ve_input(bc_pe_74_io_ve_input),
    .io_input_valid(bc_pe_74_io_input_valid),
    .io_iormac(bc_pe_74_io_iormac),
    .io_ve_out(bc_pe_74_io_ve_out),
    .io_ho_out(bc_pe_74_io_ho_out),
    .io_res_out(bc_pe_74_io_res_out)
  );
  bc_pe bc_pe_75 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_75_clock),
    .reset(bc_pe_75_reset),
    .io_ho_input(bc_pe_75_io_ho_input),
    .io_ve_input(bc_pe_75_io_ve_input),
    .io_input_valid(bc_pe_75_io_input_valid),
    .io_iormac(bc_pe_75_io_iormac),
    .io_ve_out(bc_pe_75_io_ve_out),
    .io_ho_out(bc_pe_75_io_ho_out),
    .io_res_out(bc_pe_75_io_res_out)
  );
  bc_pe bc_pe_76 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_76_clock),
    .reset(bc_pe_76_reset),
    .io_ho_input(bc_pe_76_io_ho_input),
    .io_ve_input(bc_pe_76_io_ve_input),
    .io_input_valid(bc_pe_76_io_input_valid),
    .io_iormac(bc_pe_76_io_iormac),
    .io_ve_out(bc_pe_76_io_ve_out),
    .io_ho_out(bc_pe_76_io_ho_out),
    .io_res_out(bc_pe_76_io_res_out)
  );
  bc_pe bc_pe_77 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_77_clock),
    .reset(bc_pe_77_reset),
    .io_ho_input(bc_pe_77_io_ho_input),
    .io_ve_input(bc_pe_77_io_ve_input),
    .io_input_valid(bc_pe_77_io_input_valid),
    .io_iormac(bc_pe_77_io_iormac),
    .io_ve_out(bc_pe_77_io_ve_out),
    .io_ho_out(bc_pe_77_io_ho_out),
    .io_res_out(bc_pe_77_io_res_out)
  );
  bc_pe bc_pe_78 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_78_clock),
    .reset(bc_pe_78_reset),
    .io_ho_input(bc_pe_78_io_ho_input),
    .io_ve_input(bc_pe_78_io_ve_input),
    .io_input_valid(bc_pe_78_io_input_valid),
    .io_iormac(bc_pe_78_io_iormac),
    .io_ve_out(bc_pe_78_io_ve_out),
    .io_ho_out(bc_pe_78_io_ho_out),
    .io_res_out(bc_pe_78_io_res_out)
  );
  bc_pe bc_pe_79 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_79_clock),
    .reset(bc_pe_79_reset),
    .io_ho_input(bc_pe_79_io_ho_input),
    .io_ve_input(bc_pe_79_io_ve_input),
    .io_input_valid(bc_pe_79_io_input_valid),
    .io_iormac(bc_pe_79_io_iormac),
    .io_ve_out(bc_pe_79_io_ve_out),
    .io_ho_out(bc_pe_79_io_ho_out),
    .io_res_out(bc_pe_79_io_res_out)
  );
  bc_pe bc_pe_80 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_80_clock),
    .reset(bc_pe_80_reset),
    .io_ho_input(bc_pe_80_io_ho_input),
    .io_ve_input(bc_pe_80_io_ve_input),
    .io_input_valid(bc_pe_80_io_input_valid),
    .io_iormac(bc_pe_80_io_iormac),
    .io_ve_out(bc_pe_80_io_ve_out),
    .io_ho_out(bc_pe_80_io_ho_out),
    .io_res_out(bc_pe_80_io_res_out)
  );
  bc_pe bc_pe_81 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_81_clock),
    .reset(bc_pe_81_reset),
    .io_ho_input(bc_pe_81_io_ho_input),
    .io_ve_input(bc_pe_81_io_ve_input),
    .io_input_valid(bc_pe_81_io_input_valid),
    .io_iormac(bc_pe_81_io_iormac),
    .io_ve_out(bc_pe_81_io_ve_out),
    .io_ho_out(bc_pe_81_io_ho_out),
    .io_res_out(bc_pe_81_io_res_out)
  );
  bc_pe bc_pe_82 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_82_clock),
    .reset(bc_pe_82_reset),
    .io_ho_input(bc_pe_82_io_ho_input),
    .io_ve_input(bc_pe_82_io_ve_input),
    .io_input_valid(bc_pe_82_io_input_valid),
    .io_iormac(bc_pe_82_io_iormac),
    .io_ve_out(bc_pe_82_io_ve_out),
    .io_ho_out(bc_pe_82_io_ho_out),
    .io_res_out(bc_pe_82_io_res_out)
  );
  bc_pe bc_pe_83 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_83_clock),
    .reset(bc_pe_83_reset),
    .io_ho_input(bc_pe_83_io_ho_input),
    .io_ve_input(bc_pe_83_io_ve_input),
    .io_input_valid(bc_pe_83_io_input_valid),
    .io_iormac(bc_pe_83_io_iormac),
    .io_ve_out(bc_pe_83_io_ve_out),
    .io_ho_out(bc_pe_83_io_ho_out),
    .io_res_out(bc_pe_83_io_res_out)
  );
  bc_pe bc_pe_84 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_84_clock),
    .reset(bc_pe_84_reset),
    .io_ho_input(bc_pe_84_io_ho_input),
    .io_ve_input(bc_pe_84_io_ve_input),
    .io_input_valid(bc_pe_84_io_input_valid),
    .io_iormac(bc_pe_84_io_iormac),
    .io_ve_out(bc_pe_84_io_ve_out),
    .io_ho_out(bc_pe_84_io_ho_out),
    .io_res_out(bc_pe_84_io_res_out)
  );
  bc_pe bc_pe_85 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_85_clock),
    .reset(bc_pe_85_reset),
    .io_ho_input(bc_pe_85_io_ho_input),
    .io_ve_input(bc_pe_85_io_ve_input),
    .io_input_valid(bc_pe_85_io_input_valid),
    .io_iormac(bc_pe_85_io_iormac),
    .io_ve_out(bc_pe_85_io_ve_out),
    .io_ho_out(bc_pe_85_io_ho_out),
    .io_res_out(bc_pe_85_io_res_out)
  );
  bc_pe bc_pe_86 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_86_clock),
    .reset(bc_pe_86_reset),
    .io_ho_input(bc_pe_86_io_ho_input),
    .io_ve_input(bc_pe_86_io_ve_input),
    .io_input_valid(bc_pe_86_io_input_valid),
    .io_iormac(bc_pe_86_io_iormac),
    .io_ve_out(bc_pe_86_io_ve_out),
    .io_ho_out(bc_pe_86_io_ho_out),
    .io_res_out(bc_pe_86_io_res_out)
  );
  bc_pe bc_pe_87 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_87_clock),
    .reset(bc_pe_87_reset),
    .io_ho_input(bc_pe_87_io_ho_input),
    .io_ve_input(bc_pe_87_io_ve_input),
    .io_input_valid(bc_pe_87_io_input_valid),
    .io_iormac(bc_pe_87_io_iormac),
    .io_ve_out(bc_pe_87_io_ve_out),
    .io_ho_out(bc_pe_87_io_ho_out),
    .io_res_out(bc_pe_87_io_res_out)
  );
  bc_pe bc_pe_88 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_88_clock),
    .reset(bc_pe_88_reset),
    .io_ho_input(bc_pe_88_io_ho_input),
    .io_ve_input(bc_pe_88_io_ve_input),
    .io_input_valid(bc_pe_88_io_input_valid),
    .io_iormac(bc_pe_88_io_iormac),
    .io_ve_out(bc_pe_88_io_ve_out),
    .io_ho_out(bc_pe_88_io_ho_out),
    .io_res_out(bc_pe_88_io_res_out)
  );
  bc_pe bc_pe_89 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_89_clock),
    .reset(bc_pe_89_reset),
    .io_ho_input(bc_pe_89_io_ho_input),
    .io_ve_input(bc_pe_89_io_ve_input),
    .io_input_valid(bc_pe_89_io_input_valid),
    .io_iormac(bc_pe_89_io_iormac),
    .io_ve_out(bc_pe_89_io_ve_out),
    .io_ho_out(bc_pe_89_io_ho_out),
    .io_res_out(bc_pe_89_io_res_out)
  );
  bc_pe bc_pe_90 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_90_clock),
    .reset(bc_pe_90_reset),
    .io_ho_input(bc_pe_90_io_ho_input),
    .io_ve_input(bc_pe_90_io_ve_input),
    .io_input_valid(bc_pe_90_io_input_valid),
    .io_iormac(bc_pe_90_io_iormac),
    .io_ve_out(bc_pe_90_io_ve_out),
    .io_ho_out(bc_pe_90_io_ho_out),
    .io_res_out(bc_pe_90_io_res_out)
  );
  bc_pe bc_pe_91 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_91_clock),
    .reset(bc_pe_91_reset),
    .io_ho_input(bc_pe_91_io_ho_input),
    .io_ve_input(bc_pe_91_io_ve_input),
    .io_input_valid(bc_pe_91_io_input_valid),
    .io_iormac(bc_pe_91_io_iormac),
    .io_ve_out(bc_pe_91_io_ve_out),
    .io_ho_out(bc_pe_91_io_ho_out),
    .io_res_out(bc_pe_91_io_res_out)
  );
  bc_pe bc_pe_92 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_92_clock),
    .reset(bc_pe_92_reset),
    .io_ho_input(bc_pe_92_io_ho_input),
    .io_ve_input(bc_pe_92_io_ve_input),
    .io_input_valid(bc_pe_92_io_input_valid),
    .io_iormac(bc_pe_92_io_iormac),
    .io_ve_out(bc_pe_92_io_ve_out),
    .io_ho_out(bc_pe_92_io_ho_out),
    .io_res_out(bc_pe_92_io_res_out)
  );
  bc_pe bc_pe_93 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_93_clock),
    .reset(bc_pe_93_reset),
    .io_ho_input(bc_pe_93_io_ho_input),
    .io_ve_input(bc_pe_93_io_ve_input),
    .io_input_valid(bc_pe_93_io_input_valid),
    .io_iormac(bc_pe_93_io_iormac),
    .io_ve_out(bc_pe_93_io_ve_out),
    .io_ho_out(bc_pe_93_io_ho_out),
    .io_res_out(bc_pe_93_io_res_out)
  );
  bc_pe bc_pe_94 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_94_clock),
    .reset(bc_pe_94_reset),
    .io_ho_input(bc_pe_94_io_ho_input),
    .io_ve_input(bc_pe_94_io_ve_input),
    .io_input_valid(bc_pe_94_io_input_valid),
    .io_iormac(bc_pe_94_io_iormac),
    .io_ve_out(bc_pe_94_io_ve_out),
    .io_ho_out(bc_pe_94_io_ho_out),
    .io_res_out(bc_pe_94_io_res_out)
  );
  bc_pe bc_pe_95 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_95_clock),
    .reset(bc_pe_95_reset),
    .io_ho_input(bc_pe_95_io_ho_input),
    .io_ve_input(bc_pe_95_io_ve_input),
    .io_input_valid(bc_pe_95_io_input_valid),
    .io_iormac(bc_pe_95_io_iormac),
    .io_ve_out(bc_pe_95_io_ve_out),
    .io_ho_out(bc_pe_95_io_ho_out),
    .io_res_out(bc_pe_95_io_res_out)
  );
  bc_pe bc_pe_96 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_96_clock),
    .reset(bc_pe_96_reset),
    .io_ho_input(bc_pe_96_io_ho_input),
    .io_ve_input(bc_pe_96_io_ve_input),
    .io_input_valid(bc_pe_96_io_input_valid),
    .io_iormac(bc_pe_96_io_iormac),
    .io_ve_out(bc_pe_96_io_ve_out),
    .io_ho_out(bc_pe_96_io_ho_out),
    .io_res_out(bc_pe_96_io_res_out)
  );
  bc_pe bc_pe_97 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_97_clock),
    .reset(bc_pe_97_reset),
    .io_ho_input(bc_pe_97_io_ho_input),
    .io_ve_input(bc_pe_97_io_ve_input),
    .io_input_valid(bc_pe_97_io_input_valid),
    .io_iormac(bc_pe_97_io_iormac),
    .io_ve_out(bc_pe_97_io_ve_out),
    .io_ho_out(bc_pe_97_io_ho_out),
    .io_res_out(bc_pe_97_io_res_out)
  );
  bc_pe bc_pe_98 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_98_clock),
    .reset(bc_pe_98_reset),
    .io_ho_input(bc_pe_98_io_ho_input),
    .io_ve_input(bc_pe_98_io_ve_input),
    .io_input_valid(bc_pe_98_io_input_valid),
    .io_iormac(bc_pe_98_io_iormac),
    .io_ve_out(bc_pe_98_io_ve_out),
    .io_ho_out(bc_pe_98_io_ho_out),
    .io_res_out(bc_pe_98_io_res_out)
  );
  bc_pe bc_pe_99 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_99_clock),
    .reset(bc_pe_99_reset),
    .io_ho_input(bc_pe_99_io_ho_input),
    .io_ve_input(bc_pe_99_io_ve_input),
    .io_input_valid(bc_pe_99_io_input_valid),
    .io_iormac(bc_pe_99_io_iormac),
    .io_ve_out(bc_pe_99_io_ve_out),
    .io_ho_out(bc_pe_99_io_ho_out),
    .io_res_out(bc_pe_99_io_res_out)
  );
  bc_pe bc_pe_100 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_100_clock),
    .reset(bc_pe_100_reset),
    .io_ho_input(bc_pe_100_io_ho_input),
    .io_ve_input(bc_pe_100_io_ve_input),
    .io_input_valid(bc_pe_100_io_input_valid),
    .io_iormac(bc_pe_100_io_iormac),
    .io_ve_out(bc_pe_100_io_ve_out),
    .io_ho_out(bc_pe_100_io_ho_out),
    .io_res_out(bc_pe_100_io_res_out)
  );
  bc_pe bc_pe_101 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_101_clock),
    .reset(bc_pe_101_reset),
    .io_ho_input(bc_pe_101_io_ho_input),
    .io_ve_input(bc_pe_101_io_ve_input),
    .io_input_valid(bc_pe_101_io_input_valid),
    .io_iormac(bc_pe_101_io_iormac),
    .io_ve_out(bc_pe_101_io_ve_out),
    .io_ho_out(bc_pe_101_io_ho_out),
    .io_res_out(bc_pe_101_io_res_out)
  );
  bc_pe bc_pe_102 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_102_clock),
    .reset(bc_pe_102_reset),
    .io_ho_input(bc_pe_102_io_ho_input),
    .io_ve_input(bc_pe_102_io_ve_input),
    .io_input_valid(bc_pe_102_io_input_valid),
    .io_iormac(bc_pe_102_io_iormac),
    .io_ve_out(bc_pe_102_io_ve_out),
    .io_ho_out(bc_pe_102_io_ho_out),
    .io_res_out(bc_pe_102_io_res_out)
  );
  bc_pe bc_pe_103 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_103_clock),
    .reset(bc_pe_103_reset),
    .io_ho_input(bc_pe_103_io_ho_input),
    .io_ve_input(bc_pe_103_io_ve_input),
    .io_input_valid(bc_pe_103_io_input_valid),
    .io_iormac(bc_pe_103_io_iormac),
    .io_ve_out(bc_pe_103_io_ve_out),
    .io_ho_out(bc_pe_103_io_ho_out),
    .io_res_out(bc_pe_103_io_res_out)
  );
  bc_pe bc_pe_104 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_104_clock),
    .reset(bc_pe_104_reset),
    .io_ho_input(bc_pe_104_io_ho_input),
    .io_ve_input(bc_pe_104_io_ve_input),
    .io_input_valid(bc_pe_104_io_input_valid),
    .io_iormac(bc_pe_104_io_iormac),
    .io_ve_out(bc_pe_104_io_ve_out),
    .io_ho_out(bc_pe_104_io_ho_out),
    .io_res_out(bc_pe_104_io_res_out)
  );
  bc_pe bc_pe_105 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_105_clock),
    .reset(bc_pe_105_reset),
    .io_ho_input(bc_pe_105_io_ho_input),
    .io_ve_input(bc_pe_105_io_ve_input),
    .io_input_valid(bc_pe_105_io_input_valid),
    .io_iormac(bc_pe_105_io_iormac),
    .io_ve_out(bc_pe_105_io_ve_out),
    .io_ho_out(bc_pe_105_io_ho_out),
    .io_res_out(bc_pe_105_io_res_out)
  );
  bc_pe bc_pe_106 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_106_clock),
    .reset(bc_pe_106_reset),
    .io_ho_input(bc_pe_106_io_ho_input),
    .io_ve_input(bc_pe_106_io_ve_input),
    .io_input_valid(bc_pe_106_io_input_valid),
    .io_iormac(bc_pe_106_io_iormac),
    .io_ve_out(bc_pe_106_io_ve_out),
    .io_ho_out(bc_pe_106_io_ho_out),
    .io_res_out(bc_pe_106_io_res_out)
  );
  bc_pe bc_pe_107 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_107_clock),
    .reset(bc_pe_107_reset),
    .io_ho_input(bc_pe_107_io_ho_input),
    .io_ve_input(bc_pe_107_io_ve_input),
    .io_input_valid(bc_pe_107_io_input_valid),
    .io_iormac(bc_pe_107_io_iormac),
    .io_ve_out(bc_pe_107_io_ve_out),
    .io_ho_out(bc_pe_107_io_ho_out),
    .io_res_out(bc_pe_107_io_res_out)
  );
  bc_pe bc_pe_108 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_108_clock),
    .reset(bc_pe_108_reset),
    .io_ho_input(bc_pe_108_io_ho_input),
    .io_ve_input(bc_pe_108_io_ve_input),
    .io_input_valid(bc_pe_108_io_input_valid),
    .io_iormac(bc_pe_108_io_iormac),
    .io_ve_out(bc_pe_108_io_ve_out),
    .io_ho_out(bc_pe_108_io_ho_out),
    .io_res_out(bc_pe_108_io_res_out)
  );
  bc_pe bc_pe_109 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_109_clock),
    .reset(bc_pe_109_reset),
    .io_ho_input(bc_pe_109_io_ho_input),
    .io_ve_input(bc_pe_109_io_ve_input),
    .io_input_valid(bc_pe_109_io_input_valid),
    .io_iormac(bc_pe_109_io_iormac),
    .io_ve_out(bc_pe_109_io_ve_out),
    .io_ho_out(bc_pe_109_io_ho_out),
    .io_res_out(bc_pe_109_io_res_out)
  );
  bc_pe bc_pe_110 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_110_clock),
    .reset(bc_pe_110_reset),
    .io_ho_input(bc_pe_110_io_ho_input),
    .io_ve_input(bc_pe_110_io_ve_input),
    .io_input_valid(bc_pe_110_io_input_valid),
    .io_iormac(bc_pe_110_io_iormac),
    .io_ve_out(bc_pe_110_io_ve_out),
    .io_ho_out(bc_pe_110_io_ho_out),
    .io_res_out(bc_pe_110_io_res_out)
  );
  bc_pe bc_pe_111 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_111_clock),
    .reset(bc_pe_111_reset),
    .io_ho_input(bc_pe_111_io_ho_input),
    .io_ve_input(bc_pe_111_io_ve_input),
    .io_input_valid(bc_pe_111_io_input_valid),
    .io_iormac(bc_pe_111_io_iormac),
    .io_ve_out(bc_pe_111_io_ve_out),
    .io_ho_out(bc_pe_111_io_ho_out),
    .io_res_out(bc_pe_111_io_res_out)
  );
  bc_pe bc_pe_112 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_112_clock),
    .reset(bc_pe_112_reset),
    .io_ho_input(bc_pe_112_io_ho_input),
    .io_ve_input(bc_pe_112_io_ve_input),
    .io_input_valid(bc_pe_112_io_input_valid),
    .io_iormac(bc_pe_112_io_iormac),
    .io_ve_out(bc_pe_112_io_ve_out),
    .io_ho_out(bc_pe_112_io_ho_out),
    .io_res_out(bc_pe_112_io_res_out)
  );
  bc_pe bc_pe_113 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_113_clock),
    .reset(bc_pe_113_reset),
    .io_ho_input(bc_pe_113_io_ho_input),
    .io_ve_input(bc_pe_113_io_ve_input),
    .io_input_valid(bc_pe_113_io_input_valid),
    .io_iormac(bc_pe_113_io_iormac),
    .io_ve_out(bc_pe_113_io_ve_out),
    .io_ho_out(bc_pe_113_io_ho_out),
    .io_res_out(bc_pe_113_io_res_out)
  );
  bc_pe bc_pe_114 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_114_clock),
    .reset(bc_pe_114_reset),
    .io_ho_input(bc_pe_114_io_ho_input),
    .io_ve_input(bc_pe_114_io_ve_input),
    .io_input_valid(bc_pe_114_io_input_valid),
    .io_iormac(bc_pe_114_io_iormac),
    .io_ve_out(bc_pe_114_io_ve_out),
    .io_ho_out(bc_pe_114_io_ho_out),
    .io_res_out(bc_pe_114_io_res_out)
  );
  bc_pe bc_pe_115 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_115_clock),
    .reset(bc_pe_115_reset),
    .io_ho_input(bc_pe_115_io_ho_input),
    .io_ve_input(bc_pe_115_io_ve_input),
    .io_input_valid(bc_pe_115_io_input_valid),
    .io_iormac(bc_pe_115_io_iormac),
    .io_ve_out(bc_pe_115_io_ve_out),
    .io_ho_out(bc_pe_115_io_ho_out),
    .io_res_out(bc_pe_115_io_res_out)
  );
  bc_pe bc_pe_116 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_116_clock),
    .reset(bc_pe_116_reset),
    .io_ho_input(bc_pe_116_io_ho_input),
    .io_ve_input(bc_pe_116_io_ve_input),
    .io_input_valid(bc_pe_116_io_input_valid),
    .io_iormac(bc_pe_116_io_iormac),
    .io_ve_out(bc_pe_116_io_ve_out),
    .io_ho_out(bc_pe_116_io_ho_out),
    .io_res_out(bc_pe_116_io_res_out)
  );
  bc_pe bc_pe_117 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_117_clock),
    .reset(bc_pe_117_reset),
    .io_ho_input(bc_pe_117_io_ho_input),
    .io_ve_input(bc_pe_117_io_ve_input),
    .io_input_valid(bc_pe_117_io_input_valid),
    .io_iormac(bc_pe_117_io_iormac),
    .io_ve_out(bc_pe_117_io_ve_out),
    .io_ho_out(bc_pe_117_io_ho_out),
    .io_res_out(bc_pe_117_io_res_out)
  );
  bc_pe bc_pe_118 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_118_clock),
    .reset(bc_pe_118_reset),
    .io_ho_input(bc_pe_118_io_ho_input),
    .io_ve_input(bc_pe_118_io_ve_input),
    .io_input_valid(bc_pe_118_io_input_valid),
    .io_iormac(bc_pe_118_io_iormac),
    .io_ve_out(bc_pe_118_io_ve_out),
    .io_ho_out(bc_pe_118_io_ho_out),
    .io_res_out(bc_pe_118_io_res_out)
  );
  bc_pe bc_pe_119 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_119_clock),
    .reset(bc_pe_119_reset),
    .io_ho_input(bc_pe_119_io_ho_input),
    .io_ve_input(bc_pe_119_io_ve_input),
    .io_input_valid(bc_pe_119_io_input_valid),
    .io_iormac(bc_pe_119_io_iormac),
    .io_ve_out(bc_pe_119_io_ve_out),
    .io_ho_out(bc_pe_119_io_ho_out),
    .io_res_out(bc_pe_119_io_res_out)
  );
  bc_pe bc_pe_120 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_120_clock),
    .reset(bc_pe_120_reset),
    .io_ho_input(bc_pe_120_io_ho_input),
    .io_ve_input(bc_pe_120_io_ve_input),
    .io_input_valid(bc_pe_120_io_input_valid),
    .io_iormac(bc_pe_120_io_iormac),
    .io_ve_out(bc_pe_120_io_ve_out),
    .io_ho_out(bc_pe_120_io_ho_out),
    .io_res_out(bc_pe_120_io_res_out)
  );
  bc_pe bc_pe_121 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_121_clock),
    .reset(bc_pe_121_reset),
    .io_ho_input(bc_pe_121_io_ho_input),
    .io_ve_input(bc_pe_121_io_ve_input),
    .io_input_valid(bc_pe_121_io_input_valid),
    .io_iormac(bc_pe_121_io_iormac),
    .io_ve_out(bc_pe_121_io_ve_out),
    .io_ho_out(bc_pe_121_io_ho_out),
    .io_res_out(bc_pe_121_io_res_out)
  );
  bc_pe bc_pe_122 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_122_clock),
    .reset(bc_pe_122_reset),
    .io_ho_input(bc_pe_122_io_ho_input),
    .io_ve_input(bc_pe_122_io_ve_input),
    .io_input_valid(bc_pe_122_io_input_valid),
    .io_iormac(bc_pe_122_io_iormac),
    .io_ve_out(bc_pe_122_io_ve_out),
    .io_ho_out(bc_pe_122_io_ho_out),
    .io_res_out(bc_pe_122_io_res_out)
  );
  bc_pe bc_pe_123 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_123_clock),
    .reset(bc_pe_123_reset),
    .io_ho_input(bc_pe_123_io_ho_input),
    .io_ve_input(bc_pe_123_io_ve_input),
    .io_input_valid(bc_pe_123_io_input_valid),
    .io_iormac(bc_pe_123_io_iormac),
    .io_ve_out(bc_pe_123_io_ve_out),
    .io_ho_out(bc_pe_123_io_ho_out),
    .io_res_out(bc_pe_123_io_res_out)
  );
  bc_pe bc_pe_124 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_124_clock),
    .reset(bc_pe_124_reset),
    .io_ho_input(bc_pe_124_io_ho_input),
    .io_ve_input(bc_pe_124_io_ve_input),
    .io_input_valid(bc_pe_124_io_input_valid),
    .io_iormac(bc_pe_124_io_iormac),
    .io_ve_out(bc_pe_124_io_ve_out),
    .io_ho_out(bc_pe_124_io_ho_out),
    .io_res_out(bc_pe_124_io_res_out)
  );
  bc_pe bc_pe_125 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_125_clock),
    .reset(bc_pe_125_reset),
    .io_ho_input(bc_pe_125_io_ho_input),
    .io_ve_input(bc_pe_125_io_ve_input),
    .io_input_valid(bc_pe_125_io_input_valid),
    .io_iormac(bc_pe_125_io_iormac),
    .io_ve_out(bc_pe_125_io_ve_out),
    .io_ho_out(bc_pe_125_io_ho_out),
    .io_res_out(bc_pe_125_io_res_out)
  );
  bc_pe bc_pe_126 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_126_clock),
    .reset(bc_pe_126_reset),
    .io_ho_input(bc_pe_126_io_ho_input),
    .io_ve_input(bc_pe_126_io_ve_input),
    .io_input_valid(bc_pe_126_io_input_valid),
    .io_iormac(bc_pe_126_io_iormac),
    .io_ve_out(bc_pe_126_io_ve_out),
    .io_ho_out(bc_pe_126_io_ho_out),
    .io_res_out(bc_pe_126_io_res_out)
  );
  bc_pe bc_pe_127 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_127_clock),
    .reset(bc_pe_127_reset),
    .io_ho_input(bc_pe_127_io_ho_input),
    .io_ve_input(bc_pe_127_io_ve_input),
    .io_input_valid(bc_pe_127_io_input_valid),
    .io_iormac(bc_pe_127_io_iormac),
    .io_ve_out(bc_pe_127_io_ve_out),
    .io_ho_out(bc_pe_127_io_ho_out),
    .io_res_out(bc_pe_127_io_res_out)
  );
  bc_pe bc_pe_128 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_128_clock),
    .reset(bc_pe_128_reset),
    .io_ho_input(bc_pe_128_io_ho_input),
    .io_ve_input(bc_pe_128_io_ve_input),
    .io_input_valid(bc_pe_128_io_input_valid),
    .io_iormac(bc_pe_128_io_iormac),
    .io_ve_out(bc_pe_128_io_ve_out),
    .io_ho_out(bc_pe_128_io_ho_out),
    .io_res_out(bc_pe_128_io_res_out)
  );
  bc_pe bc_pe_129 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_129_clock),
    .reset(bc_pe_129_reset),
    .io_ho_input(bc_pe_129_io_ho_input),
    .io_ve_input(bc_pe_129_io_ve_input),
    .io_input_valid(bc_pe_129_io_input_valid),
    .io_iormac(bc_pe_129_io_iormac),
    .io_ve_out(bc_pe_129_io_ve_out),
    .io_ho_out(bc_pe_129_io_ho_out),
    .io_res_out(bc_pe_129_io_res_out)
  );
  bc_pe bc_pe_130 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_130_clock),
    .reset(bc_pe_130_reset),
    .io_ho_input(bc_pe_130_io_ho_input),
    .io_ve_input(bc_pe_130_io_ve_input),
    .io_input_valid(bc_pe_130_io_input_valid),
    .io_iormac(bc_pe_130_io_iormac),
    .io_ve_out(bc_pe_130_io_ve_out),
    .io_ho_out(bc_pe_130_io_ho_out),
    .io_res_out(bc_pe_130_io_res_out)
  );
  bc_pe bc_pe_131 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_131_clock),
    .reset(bc_pe_131_reset),
    .io_ho_input(bc_pe_131_io_ho_input),
    .io_ve_input(bc_pe_131_io_ve_input),
    .io_input_valid(bc_pe_131_io_input_valid),
    .io_iormac(bc_pe_131_io_iormac),
    .io_ve_out(bc_pe_131_io_ve_out),
    .io_ho_out(bc_pe_131_io_ho_out),
    .io_res_out(bc_pe_131_io_res_out)
  );
  bc_pe bc_pe_132 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_132_clock),
    .reset(bc_pe_132_reset),
    .io_ho_input(bc_pe_132_io_ho_input),
    .io_ve_input(bc_pe_132_io_ve_input),
    .io_input_valid(bc_pe_132_io_input_valid),
    .io_iormac(bc_pe_132_io_iormac),
    .io_ve_out(bc_pe_132_io_ve_out),
    .io_ho_out(bc_pe_132_io_ho_out),
    .io_res_out(bc_pe_132_io_res_out)
  );
  bc_pe bc_pe_133 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_133_clock),
    .reset(bc_pe_133_reset),
    .io_ho_input(bc_pe_133_io_ho_input),
    .io_ve_input(bc_pe_133_io_ve_input),
    .io_input_valid(bc_pe_133_io_input_valid),
    .io_iormac(bc_pe_133_io_iormac),
    .io_ve_out(bc_pe_133_io_ve_out),
    .io_ho_out(bc_pe_133_io_ho_out),
    .io_res_out(bc_pe_133_io_res_out)
  );
  bc_pe bc_pe_134 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_134_clock),
    .reset(bc_pe_134_reset),
    .io_ho_input(bc_pe_134_io_ho_input),
    .io_ve_input(bc_pe_134_io_ve_input),
    .io_input_valid(bc_pe_134_io_input_valid),
    .io_iormac(bc_pe_134_io_iormac),
    .io_ve_out(bc_pe_134_io_ve_out),
    .io_ho_out(bc_pe_134_io_ho_out),
    .io_res_out(bc_pe_134_io_res_out)
  );
  bc_pe bc_pe_135 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_135_clock),
    .reset(bc_pe_135_reset),
    .io_ho_input(bc_pe_135_io_ho_input),
    .io_ve_input(bc_pe_135_io_ve_input),
    .io_input_valid(bc_pe_135_io_input_valid),
    .io_iormac(bc_pe_135_io_iormac),
    .io_ve_out(bc_pe_135_io_ve_out),
    .io_ho_out(bc_pe_135_io_ho_out),
    .io_res_out(bc_pe_135_io_res_out)
  );
  bc_pe bc_pe_136 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_136_clock),
    .reset(bc_pe_136_reset),
    .io_ho_input(bc_pe_136_io_ho_input),
    .io_ve_input(bc_pe_136_io_ve_input),
    .io_input_valid(bc_pe_136_io_input_valid),
    .io_iormac(bc_pe_136_io_iormac),
    .io_ve_out(bc_pe_136_io_ve_out),
    .io_ho_out(bc_pe_136_io_ho_out),
    .io_res_out(bc_pe_136_io_res_out)
  );
  bc_pe bc_pe_137 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_137_clock),
    .reset(bc_pe_137_reset),
    .io_ho_input(bc_pe_137_io_ho_input),
    .io_ve_input(bc_pe_137_io_ve_input),
    .io_input_valid(bc_pe_137_io_input_valid),
    .io_iormac(bc_pe_137_io_iormac),
    .io_ve_out(bc_pe_137_io_ve_out),
    .io_ho_out(bc_pe_137_io_ho_out),
    .io_res_out(bc_pe_137_io_res_out)
  );
  bc_pe bc_pe_138 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_138_clock),
    .reset(bc_pe_138_reset),
    .io_ho_input(bc_pe_138_io_ho_input),
    .io_ve_input(bc_pe_138_io_ve_input),
    .io_input_valid(bc_pe_138_io_input_valid),
    .io_iormac(bc_pe_138_io_iormac),
    .io_ve_out(bc_pe_138_io_ve_out),
    .io_ho_out(bc_pe_138_io_ho_out),
    .io_res_out(bc_pe_138_io_res_out)
  );
  bc_pe bc_pe_139 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_139_clock),
    .reset(bc_pe_139_reset),
    .io_ho_input(bc_pe_139_io_ho_input),
    .io_ve_input(bc_pe_139_io_ve_input),
    .io_input_valid(bc_pe_139_io_input_valid),
    .io_iormac(bc_pe_139_io_iormac),
    .io_ve_out(bc_pe_139_io_ve_out),
    .io_ho_out(bc_pe_139_io_ho_out),
    .io_res_out(bc_pe_139_io_res_out)
  );
  bc_pe bc_pe_140 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_140_clock),
    .reset(bc_pe_140_reset),
    .io_ho_input(bc_pe_140_io_ho_input),
    .io_ve_input(bc_pe_140_io_ve_input),
    .io_input_valid(bc_pe_140_io_input_valid),
    .io_iormac(bc_pe_140_io_iormac),
    .io_ve_out(bc_pe_140_io_ve_out),
    .io_ho_out(bc_pe_140_io_ho_out),
    .io_res_out(bc_pe_140_io_res_out)
  );
  bc_pe bc_pe_141 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_141_clock),
    .reset(bc_pe_141_reset),
    .io_ho_input(bc_pe_141_io_ho_input),
    .io_ve_input(bc_pe_141_io_ve_input),
    .io_input_valid(bc_pe_141_io_input_valid),
    .io_iormac(bc_pe_141_io_iormac),
    .io_ve_out(bc_pe_141_io_ve_out),
    .io_ho_out(bc_pe_141_io_ho_out),
    .io_res_out(bc_pe_141_io_res_out)
  );
  bc_pe bc_pe_142 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_142_clock),
    .reset(bc_pe_142_reset),
    .io_ho_input(bc_pe_142_io_ho_input),
    .io_ve_input(bc_pe_142_io_ve_input),
    .io_input_valid(bc_pe_142_io_input_valid),
    .io_iormac(bc_pe_142_io_iormac),
    .io_ve_out(bc_pe_142_io_ve_out),
    .io_ho_out(bc_pe_142_io_ho_out),
    .io_res_out(bc_pe_142_io_res_out)
  );
  bc_pe bc_pe_143 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_143_clock),
    .reset(bc_pe_143_reset),
    .io_ho_input(bc_pe_143_io_ho_input),
    .io_ve_input(bc_pe_143_io_ve_input),
    .io_input_valid(bc_pe_143_io_input_valid),
    .io_iormac(bc_pe_143_io_iormac),
    .io_ve_out(bc_pe_143_io_ve_out),
    .io_ho_out(bc_pe_143_io_ho_out),
    .io_res_out(bc_pe_143_io_res_out)
  );
  bc_pe bc_pe_144 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_144_clock),
    .reset(bc_pe_144_reset),
    .io_ho_input(bc_pe_144_io_ho_input),
    .io_ve_input(bc_pe_144_io_ve_input),
    .io_input_valid(bc_pe_144_io_input_valid),
    .io_iormac(bc_pe_144_io_iormac),
    .io_ve_out(bc_pe_144_io_ve_out),
    .io_ho_out(bc_pe_144_io_ho_out),
    .io_res_out(bc_pe_144_io_res_out)
  );
  bc_pe bc_pe_145 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_145_clock),
    .reset(bc_pe_145_reset),
    .io_ho_input(bc_pe_145_io_ho_input),
    .io_ve_input(bc_pe_145_io_ve_input),
    .io_input_valid(bc_pe_145_io_input_valid),
    .io_iormac(bc_pe_145_io_iormac),
    .io_ve_out(bc_pe_145_io_ve_out),
    .io_ho_out(bc_pe_145_io_ho_out),
    .io_res_out(bc_pe_145_io_res_out)
  );
  bc_pe bc_pe_146 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_146_clock),
    .reset(bc_pe_146_reset),
    .io_ho_input(bc_pe_146_io_ho_input),
    .io_ve_input(bc_pe_146_io_ve_input),
    .io_input_valid(bc_pe_146_io_input_valid),
    .io_iormac(bc_pe_146_io_iormac),
    .io_ve_out(bc_pe_146_io_ve_out),
    .io_ho_out(bc_pe_146_io_ho_out),
    .io_res_out(bc_pe_146_io_res_out)
  );
  bc_pe bc_pe_147 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_147_clock),
    .reset(bc_pe_147_reset),
    .io_ho_input(bc_pe_147_io_ho_input),
    .io_ve_input(bc_pe_147_io_ve_input),
    .io_input_valid(bc_pe_147_io_input_valid),
    .io_iormac(bc_pe_147_io_iormac),
    .io_ve_out(bc_pe_147_io_ve_out),
    .io_ho_out(bc_pe_147_io_ho_out),
    .io_res_out(bc_pe_147_io_res_out)
  );
  bc_pe bc_pe_148 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_148_clock),
    .reset(bc_pe_148_reset),
    .io_ho_input(bc_pe_148_io_ho_input),
    .io_ve_input(bc_pe_148_io_ve_input),
    .io_input_valid(bc_pe_148_io_input_valid),
    .io_iormac(bc_pe_148_io_iormac),
    .io_ve_out(bc_pe_148_io_ve_out),
    .io_ho_out(bc_pe_148_io_ho_out),
    .io_res_out(bc_pe_148_io_res_out)
  );
  bc_pe bc_pe_149 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_149_clock),
    .reset(bc_pe_149_reset),
    .io_ho_input(bc_pe_149_io_ho_input),
    .io_ve_input(bc_pe_149_io_ve_input),
    .io_input_valid(bc_pe_149_io_input_valid),
    .io_iormac(bc_pe_149_io_iormac),
    .io_ve_out(bc_pe_149_io_ve_out),
    .io_ho_out(bc_pe_149_io_ho_out),
    .io_res_out(bc_pe_149_io_res_out)
  );
  bc_pe bc_pe_150 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_150_clock),
    .reset(bc_pe_150_reset),
    .io_ho_input(bc_pe_150_io_ho_input),
    .io_ve_input(bc_pe_150_io_ve_input),
    .io_input_valid(bc_pe_150_io_input_valid),
    .io_iormac(bc_pe_150_io_iormac),
    .io_ve_out(bc_pe_150_io_ve_out),
    .io_ho_out(bc_pe_150_io_ho_out),
    .io_res_out(bc_pe_150_io_res_out)
  );
  bc_pe bc_pe_151 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_151_clock),
    .reset(bc_pe_151_reset),
    .io_ho_input(bc_pe_151_io_ho_input),
    .io_ve_input(bc_pe_151_io_ve_input),
    .io_input_valid(bc_pe_151_io_input_valid),
    .io_iormac(bc_pe_151_io_iormac),
    .io_ve_out(bc_pe_151_io_ve_out),
    .io_ho_out(bc_pe_151_io_ho_out),
    .io_res_out(bc_pe_151_io_res_out)
  );
  bc_pe bc_pe_152 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_152_clock),
    .reset(bc_pe_152_reset),
    .io_ho_input(bc_pe_152_io_ho_input),
    .io_ve_input(bc_pe_152_io_ve_input),
    .io_input_valid(bc_pe_152_io_input_valid),
    .io_iormac(bc_pe_152_io_iormac),
    .io_ve_out(bc_pe_152_io_ve_out),
    .io_ho_out(bc_pe_152_io_ho_out),
    .io_res_out(bc_pe_152_io_res_out)
  );
  bc_pe bc_pe_153 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_153_clock),
    .reset(bc_pe_153_reset),
    .io_ho_input(bc_pe_153_io_ho_input),
    .io_ve_input(bc_pe_153_io_ve_input),
    .io_input_valid(bc_pe_153_io_input_valid),
    .io_iormac(bc_pe_153_io_iormac),
    .io_ve_out(bc_pe_153_io_ve_out),
    .io_ho_out(bc_pe_153_io_ho_out),
    .io_res_out(bc_pe_153_io_res_out)
  );
  bc_pe bc_pe_154 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_154_clock),
    .reset(bc_pe_154_reset),
    .io_ho_input(bc_pe_154_io_ho_input),
    .io_ve_input(bc_pe_154_io_ve_input),
    .io_input_valid(bc_pe_154_io_input_valid),
    .io_iormac(bc_pe_154_io_iormac),
    .io_ve_out(bc_pe_154_io_ve_out),
    .io_ho_out(bc_pe_154_io_ho_out),
    .io_res_out(bc_pe_154_io_res_out)
  );
  bc_pe bc_pe_155 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_155_clock),
    .reset(bc_pe_155_reset),
    .io_ho_input(bc_pe_155_io_ho_input),
    .io_ve_input(bc_pe_155_io_ve_input),
    .io_input_valid(bc_pe_155_io_input_valid),
    .io_iormac(bc_pe_155_io_iormac),
    .io_ve_out(bc_pe_155_io_ve_out),
    .io_ho_out(bc_pe_155_io_ho_out),
    .io_res_out(bc_pe_155_io_res_out)
  );
  bc_pe bc_pe_156 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_156_clock),
    .reset(bc_pe_156_reset),
    .io_ho_input(bc_pe_156_io_ho_input),
    .io_ve_input(bc_pe_156_io_ve_input),
    .io_input_valid(bc_pe_156_io_input_valid),
    .io_iormac(bc_pe_156_io_iormac),
    .io_ve_out(bc_pe_156_io_ve_out),
    .io_ho_out(bc_pe_156_io_ho_out),
    .io_res_out(bc_pe_156_io_res_out)
  );
  bc_pe bc_pe_157 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_157_clock),
    .reset(bc_pe_157_reset),
    .io_ho_input(bc_pe_157_io_ho_input),
    .io_ve_input(bc_pe_157_io_ve_input),
    .io_input_valid(bc_pe_157_io_input_valid),
    .io_iormac(bc_pe_157_io_iormac),
    .io_ve_out(bc_pe_157_io_ve_out),
    .io_ho_out(bc_pe_157_io_ho_out),
    .io_res_out(bc_pe_157_io_res_out)
  );
  bc_pe bc_pe_158 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_158_clock),
    .reset(bc_pe_158_reset),
    .io_ho_input(bc_pe_158_io_ho_input),
    .io_ve_input(bc_pe_158_io_ve_input),
    .io_input_valid(bc_pe_158_io_input_valid),
    .io_iormac(bc_pe_158_io_iormac),
    .io_ve_out(bc_pe_158_io_ve_out),
    .io_ho_out(bc_pe_158_io_ho_out),
    .io_res_out(bc_pe_158_io_res_out)
  );
  bc_pe bc_pe_159 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_159_clock),
    .reset(bc_pe_159_reset),
    .io_ho_input(bc_pe_159_io_ho_input),
    .io_ve_input(bc_pe_159_io_ve_input),
    .io_input_valid(bc_pe_159_io_input_valid),
    .io_iormac(bc_pe_159_io_iormac),
    .io_ve_out(bc_pe_159_io_ve_out),
    .io_ho_out(bc_pe_159_io_ho_out),
    .io_res_out(bc_pe_159_io_res_out)
  );
  bc_pe bc_pe_160 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_160_clock),
    .reset(bc_pe_160_reset),
    .io_ho_input(bc_pe_160_io_ho_input),
    .io_ve_input(bc_pe_160_io_ve_input),
    .io_input_valid(bc_pe_160_io_input_valid),
    .io_iormac(bc_pe_160_io_iormac),
    .io_ve_out(bc_pe_160_io_ve_out),
    .io_ho_out(bc_pe_160_io_ho_out),
    .io_res_out(bc_pe_160_io_res_out)
  );
  bc_pe bc_pe_161 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_161_clock),
    .reset(bc_pe_161_reset),
    .io_ho_input(bc_pe_161_io_ho_input),
    .io_ve_input(bc_pe_161_io_ve_input),
    .io_input_valid(bc_pe_161_io_input_valid),
    .io_iormac(bc_pe_161_io_iormac),
    .io_ve_out(bc_pe_161_io_ve_out),
    .io_ho_out(bc_pe_161_io_ho_out),
    .io_res_out(bc_pe_161_io_res_out)
  );
  bc_pe bc_pe_162 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_162_clock),
    .reset(bc_pe_162_reset),
    .io_ho_input(bc_pe_162_io_ho_input),
    .io_ve_input(bc_pe_162_io_ve_input),
    .io_input_valid(bc_pe_162_io_input_valid),
    .io_iormac(bc_pe_162_io_iormac),
    .io_ve_out(bc_pe_162_io_ve_out),
    .io_ho_out(bc_pe_162_io_ho_out),
    .io_res_out(bc_pe_162_io_res_out)
  );
  bc_pe bc_pe_163 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_163_clock),
    .reset(bc_pe_163_reset),
    .io_ho_input(bc_pe_163_io_ho_input),
    .io_ve_input(bc_pe_163_io_ve_input),
    .io_input_valid(bc_pe_163_io_input_valid),
    .io_iormac(bc_pe_163_io_iormac),
    .io_ve_out(bc_pe_163_io_ve_out),
    .io_ho_out(bc_pe_163_io_ho_out),
    .io_res_out(bc_pe_163_io_res_out)
  );
  bc_pe bc_pe_164 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_164_clock),
    .reset(bc_pe_164_reset),
    .io_ho_input(bc_pe_164_io_ho_input),
    .io_ve_input(bc_pe_164_io_ve_input),
    .io_input_valid(bc_pe_164_io_input_valid),
    .io_iormac(bc_pe_164_io_iormac),
    .io_ve_out(bc_pe_164_io_ve_out),
    .io_ho_out(bc_pe_164_io_ho_out),
    .io_res_out(bc_pe_164_io_res_out)
  );
  bc_pe bc_pe_165 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_165_clock),
    .reset(bc_pe_165_reset),
    .io_ho_input(bc_pe_165_io_ho_input),
    .io_ve_input(bc_pe_165_io_ve_input),
    .io_input_valid(bc_pe_165_io_input_valid),
    .io_iormac(bc_pe_165_io_iormac),
    .io_ve_out(bc_pe_165_io_ve_out),
    .io_ho_out(bc_pe_165_io_ho_out),
    .io_res_out(bc_pe_165_io_res_out)
  );
  bc_pe bc_pe_166 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_166_clock),
    .reset(bc_pe_166_reset),
    .io_ho_input(bc_pe_166_io_ho_input),
    .io_ve_input(bc_pe_166_io_ve_input),
    .io_input_valid(bc_pe_166_io_input_valid),
    .io_iormac(bc_pe_166_io_iormac),
    .io_ve_out(bc_pe_166_io_ve_out),
    .io_ho_out(bc_pe_166_io_ho_out),
    .io_res_out(bc_pe_166_io_res_out)
  );
  bc_pe bc_pe_167 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_167_clock),
    .reset(bc_pe_167_reset),
    .io_ho_input(bc_pe_167_io_ho_input),
    .io_ve_input(bc_pe_167_io_ve_input),
    .io_input_valid(bc_pe_167_io_input_valid),
    .io_iormac(bc_pe_167_io_iormac),
    .io_ve_out(bc_pe_167_io_ve_out),
    .io_ho_out(bc_pe_167_io_ho_out),
    .io_res_out(bc_pe_167_io_res_out)
  );
  bc_pe bc_pe_168 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_168_clock),
    .reset(bc_pe_168_reset),
    .io_ho_input(bc_pe_168_io_ho_input),
    .io_ve_input(bc_pe_168_io_ve_input),
    .io_input_valid(bc_pe_168_io_input_valid),
    .io_iormac(bc_pe_168_io_iormac),
    .io_ve_out(bc_pe_168_io_ve_out),
    .io_ho_out(bc_pe_168_io_ho_out),
    .io_res_out(bc_pe_168_io_res_out)
  );
  bc_pe bc_pe_169 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_169_clock),
    .reset(bc_pe_169_reset),
    .io_ho_input(bc_pe_169_io_ho_input),
    .io_ve_input(bc_pe_169_io_ve_input),
    .io_input_valid(bc_pe_169_io_input_valid),
    .io_iormac(bc_pe_169_io_iormac),
    .io_ve_out(bc_pe_169_io_ve_out),
    .io_ho_out(bc_pe_169_io_ho_out),
    .io_res_out(bc_pe_169_io_res_out)
  );
  bc_pe bc_pe_170 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_170_clock),
    .reset(bc_pe_170_reset),
    .io_ho_input(bc_pe_170_io_ho_input),
    .io_ve_input(bc_pe_170_io_ve_input),
    .io_input_valid(bc_pe_170_io_input_valid),
    .io_iormac(bc_pe_170_io_iormac),
    .io_ve_out(bc_pe_170_io_ve_out),
    .io_ho_out(bc_pe_170_io_ho_out),
    .io_res_out(bc_pe_170_io_res_out)
  );
  bc_pe bc_pe_171 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_171_clock),
    .reset(bc_pe_171_reset),
    .io_ho_input(bc_pe_171_io_ho_input),
    .io_ve_input(bc_pe_171_io_ve_input),
    .io_input_valid(bc_pe_171_io_input_valid),
    .io_iormac(bc_pe_171_io_iormac),
    .io_ve_out(bc_pe_171_io_ve_out),
    .io_ho_out(bc_pe_171_io_ho_out),
    .io_res_out(bc_pe_171_io_res_out)
  );
  bc_pe bc_pe_172 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_172_clock),
    .reset(bc_pe_172_reset),
    .io_ho_input(bc_pe_172_io_ho_input),
    .io_ve_input(bc_pe_172_io_ve_input),
    .io_input_valid(bc_pe_172_io_input_valid),
    .io_iormac(bc_pe_172_io_iormac),
    .io_ve_out(bc_pe_172_io_ve_out),
    .io_ho_out(bc_pe_172_io_ho_out),
    .io_res_out(bc_pe_172_io_res_out)
  );
  bc_pe bc_pe_173 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_173_clock),
    .reset(bc_pe_173_reset),
    .io_ho_input(bc_pe_173_io_ho_input),
    .io_ve_input(bc_pe_173_io_ve_input),
    .io_input_valid(bc_pe_173_io_input_valid),
    .io_iormac(bc_pe_173_io_iormac),
    .io_ve_out(bc_pe_173_io_ve_out),
    .io_ho_out(bc_pe_173_io_ho_out),
    .io_res_out(bc_pe_173_io_res_out)
  );
  bc_pe bc_pe_174 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_174_clock),
    .reset(bc_pe_174_reset),
    .io_ho_input(bc_pe_174_io_ho_input),
    .io_ve_input(bc_pe_174_io_ve_input),
    .io_input_valid(bc_pe_174_io_input_valid),
    .io_iormac(bc_pe_174_io_iormac),
    .io_ve_out(bc_pe_174_io_ve_out),
    .io_ho_out(bc_pe_174_io_ho_out),
    .io_res_out(bc_pe_174_io_res_out)
  );
  bc_pe bc_pe_175 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_175_clock),
    .reset(bc_pe_175_reset),
    .io_ho_input(bc_pe_175_io_ho_input),
    .io_ve_input(bc_pe_175_io_ve_input),
    .io_input_valid(bc_pe_175_io_input_valid),
    .io_iormac(bc_pe_175_io_iormac),
    .io_ve_out(bc_pe_175_io_ve_out),
    .io_ho_out(bc_pe_175_io_ho_out),
    .io_res_out(bc_pe_175_io_res_out)
  );
  bc_pe bc_pe_176 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_176_clock),
    .reset(bc_pe_176_reset),
    .io_ho_input(bc_pe_176_io_ho_input),
    .io_ve_input(bc_pe_176_io_ve_input),
    .io_input_valid(bc_pe_176_io_input_valid),
    .io_iormac(bc_pe_176_io_iormac),
    .io_ve_out(bc_pe_176_io_ve_out),
    .io_ho_out(bc_pe_176_io_ho_out),
    .io_res_out(bc_pe_176_io_res_out)
  );
  bc_pe bc_pe_177 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_177_clock),
    .reset(bc_pe_177_reset),
    .io_ho_input(bc_pe_177_io_ho_input),
    .io_ve_input(bc_pe_177_io_ve_input),
    .io_input_valid(bc_pe_177_io_input_valid),
    .io_iormac(bc_pe_177_io_iormac),
    .io_ve_out(bc_pe_177_io_ve_out),
    .io_ho_out(bc_pe_177_io_ho_out),
    .io_res_out(bc_pe_177_io_res_out)
  );
  bc_pe bc_pe_178 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_178_clock),
    .reset(bc_pe_178_reset),
    .io_ho_input(bc_pe_178_io_ho_input),
    .io_ve_input(bc_pe_178_io_ve_input),
    .io_input_valid(bc_pe_178_io_input_valid),
    .io_iormac(bc_pe_178_io_iormac),
    .io_ve_out(bc_pe_178_io_ve_out),
    .io_ho_out(bc_pe_178_io_ho_out),
    .io_res_out(bc_pe_178_io_res_out)
  );
  bc_pe bc_pe_179 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_179_clock),
    .reset(bc_pe_179_reset),
    .io_ho_input(bc_pe_179_io_ho_input),
    .io_ve_input(bc_pe_179_io_ve_input),
    .io_input_valid(bc_pe_179_io_input_valid),
    .io_iormac(bc_pe_179_io_iormac),
    .io_ve_out(bc_pe_179_io_ve_out),
    .io_ho_out(bc_pe_179_io_ho_out),
    .io_res_out(bc_pe_179_io_res_out)
  );
  bc_pe bc_pe_180 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_180_clock),
    .reset(bc_pe_180_reset),
    .io_ho_input(bc_pe_180_io_ho_input),
    .io_ve_input(bc_pe_180_io_ve_input),
    .io_input_valid(bc_pe_180_io_input_valid),
    .io_iormac(bc_pe_180_io_iormac),
    .io_ve_out(bc_pe_180_io_ve_out),
    .io_ho_out(bc_pe_180_io_ho_out),
    .io_res_out(bc_pe_180_io_res_out)
  );
  bc_pe bc_pe_181 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_181_clock),
    .reset(bc_pe_181_reset),
    .io_ho_input(bc_pe_181_io_ho_input),
    .io_ve_input(bc_pe_181_io_ve_input),
    .io_input_valid(bc_pe_181_io_input_valid),
    .io_iormac(bc_pe_181_io_iormac),
    .io_ve_out(bc_pe_181_io_ve_out),
    .io_ho_out(bc_pe_181_io_ho_out),
    .io_res_out(bc_pe_181_io_res_out)
  );
  bc_pe bc_pe_182 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_182_clock),
    .reset(bc_pe_182_reset),
    .io_ho_input(bc_pe_182_io_ho_input),
    .io_ve_input(bc_pe_182_io_ve_input),
    .io_input_valid(bc_pe_182_io_input_valid),
    .io_iormac(bc_pe_182_io_iormac),
    .io_ve_out(bc_pe_182_io_ve_out),
    .io_ho_out(bc_pe_182_io_ho_out),
    .io_res_out(bc_pe_182_io_res_out)
  );
  bc_pe bc_pe_183 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_183_clock),
    .reset(bc_pe_183_reset),
    .io_ho_input(bc_pe_183_io_ho_input),
    .io_ve_input(bc_pe_183_io_ve_input),
    .io_input_valid(bc_pe_183_io_input_valid),
    .io_iormac(bc_pe_183_io_iormac),
    .io_ve_out(bc_pe_183_io_ve_out),
    .io_ho_out(bc_pe_183_io_ho_out),
    .io_res_out(bc_pe_183_io_res_out)
  );
  bc_pe bc_pe_184 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_184_clock),
    .reset(bc_pe_184_reset),
    .io_ho_input(bc_pe_184_io_ho_input),
    .io_ve_input(bc_pe_184_io_ve_input),
    .io_input_valid(bc_pe_184_io_input_valid),
    .io_iormac(bc_pe_184_io_iormac),
    .io_ve_out(bc_pe_184_io_ve_out),
    .io_ho_out(bc_pe_184_io_ho_out),
    .io_res_out(bc_pe_184_io_res_out)
  );
  bc_pe bc_pe_185 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_185_clock),
    .reset(bc_pe_185_reset),
    .io_ho_input(bc_pe_185_io_ho_input),
    .io_ve_input(bc_pe_185_io_ve_input),
    .io_input_valid(bc_pe_185_io_input_valid),
    .io_iormac(bc_pe_185_io_iormac),
    .io_ve_out(bc_pe_185_io_ve_out),
    .io_ho_out(bc_pe_185_io_ho_out),
    .io_res_out(bc_pe_185_io_res_out)
  );
  bc_pe bc_pe_186 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_186_clock),
    .reset(bc_pe_186_reset),
    .io_ho_input(bc_pe_186_io_ho_input),
    .io_ve_input(bc_pe_186_io_ve_input),
    .io_input_valid(bc_pe_186_io_input_valid),
    .io_iormac(bc_pe_186_io_iormac),
    .io_ve_out(bc_pe_186_io_ve_out),
    .io_ho_out(bc_pe_186_io_ho_out),
    .io_res_out(bc_pe_186_io_res_out)
  );
  bc_pe bc_pe_187 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_187_clock),
    .reset(bc_pe_187_reset),
    .io_ho_input(bc_pe_187_io_ho_input),
    .io_ve_input(bc_pe_187_io_ve_input),
    .io_input_valid(bc_pe_187_io_input_valid),
    .io_iormac(bc_pe_187_io_iormac),
    .io_ve_out(bc_pe_187_io_ve_out),
    .io_ho_out(bc_pe_187_io_ho_out),
    .io_res_out(bc_pe_187_io_res_out)
  );
  bc_pe bc_pe_188 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_188_clock),
    .reset(bc_pe_188_reset),
    .io_ho_input(bc_pe_188_io_ho_input),
    .io_ve_input(bc_pe_188_io_ve_input),
    .io_input_valid(bc_pe_188_io_input_valid),
    .io_iormac(bc_pe_188_io_iormac),
    .io_ve_out(bc_pe_188_io_ve_out),
    .io_ho_out(bc_pe_188_io_ho_out),
    .io_res_out(bc_pe_188_io_res_out)
  );
  bc_pe bc_pe_189 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_189_clock),
    .reset(bc_pe_189_reset),
    .io_ho_input(bc_pe_189_io_ho_input),
    .io_ve_input(bc_pe_189_io_ve_input),
    .io_input_valid(bc_pe_189_io_input_valid),
    .io_iormac(bc_pe_189_io_iormac),
    .io_ve_out(bc_pe_189_io_ve_out),
    .io_ho_out(bc_pe_189_io_ho_out),
    .io_res_out(bc_pe_189_io_res_out)
  );
  bc_pe bc_pe_190 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_190_clock),
    .reset(bc_pe_190_reset),
    .io_ho_input(bc_pe_190_io_ho_input),
    .io_ve_input(bc_pe_190_io_ve_input),
    .io_input_valid(bc_pe_190_io_input_valid),
    .io_iormac(bc_pe_190_io_iormac),
    .io_ve_out(bc_pe_190_io_ve_out),
    .io_ho_out(bc_pe_190_io_ho_out),
    .io_res_out(bc_pe_190_io_res_out)
  );
  bc_pe bc_pe_191 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_191_clock),
    .reset(bc_pe_191_reset),
    .io_ho_input(bc_pe_191_io_ho_input),
    .io_ve_input(bc_pe_191_io_ve_input),
    .io_input_valid(bc_pe_191_io_input_valid),
    .io_iormac(bc_pe_191_io_iormac),
    .io_ve_out(bc_pe_191_io_ve_out),
    .io_ho_out(bc_pe_191_io_ho_out),
    .io_res_out(bc_pe_191_io_res_out)
  );
  bc_pe bc_pe_192 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_192_clock),
    .reset(bc_pe_192_reset),
    .io_ho_input(bc_pe_192_io_ho_input),
    .io_ve_input(bc_pe_192_io_ve_input),
    .io_input_valid(bc_pe_192_io_input_valid),
    .io_iormac(bc_pe_192_io_iormac),
    .io_ve_out(bc_pe_192_io_ve_out),
    .io_ho_out(bc_pe_192_io_ho_out),
    .io_res_out(bc_pe_192_io_res_out)
  );
  bc_pe bc_pe_193 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_193_clock),
    .reset(bc_pe_193_reset),
    .io_ho_input(bc_pe_193_io_ho_input),
    .io_ve_input(bc_pe_193_io_ve_input),
    .io_input_valid(bc_pe_193_io_input_valid),
    .io_iormac(bc_pe_193_io_iormac),
    .io_ve_out(bc_pe_193_io_ve_out),
    .io_ho_out(bc_pe_193_io_ho_out),
    .io_res_out(bc_pe_193_io_res_out)
  );
  bc_pe bc_pe_194 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_194_clock),
    .reset(bc_pe_194_reset),
    .io_ho_input(bc_pe_194_io_ho_input),
    .io_ve_input(bc_pe_194_io_ve_input),
    .io_input_valid(bc_pe_194_io_input_valid),
    .io_iormac(bc_pe_194_io_iormac),
    .io_ve_out(bc_pe_194_io_ve_out),
    .io_ho_out(bc_pe_194_io_ho_out),
    .io_res_out(bc_pe_194_io_res_out)
  );
  bc_pe bc_pe_195 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_195_clock),
    .reset(bc_pe_195_reset),
    .io_ho_input(bc_pe_195_io_ho_input),
    .io_ve_input(bc_pe_195_io_ve_input),
    .io_input_valid(bc_pe_195_io_input_valid),
    .io_iormac(bc_pe_195_io_iormac),
    .io_ve_out(bc_pe_195_io_ve_out),
    .io_ho_out(bc_pe_195_io_ho_out),
    .io_res_out(bc_pe_195_io_res_out)
  );
  bc_pe bc_pe_196 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_196_clock),
    .reset(bc_pe_196_reset),
    .io_ho_input(bc_pe_196_io_ho_input),
    .io_ve_input(bc_pe_196_io_ve_input),
    .io_input_valid(bc_pe_196_io_input_valid),
    .io_iormac(bc_pe_196_io_iormac),
    .io_ve_out(bc_pe_196_io_ve_out),
    .io_ho_out(bc_pe_196_io_ho_out),
    .io_res_out(bc_pe_196_io_res_out)
  );
  bc_pe bc_pe_197 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_197_clock),
    .reset(bc_pe_197_reset),
    .io_ho_input(bc_pe_197_io_ho_input),
    .io_ve_input(bc_pe_197_io_ve_input),
    .io_input_valid(bc_pe_197_io_input_valid),
    .io_iormac(bc_pe_197_io_iormac),
    .io_ve_out(bc_pe_197_io_ve_out),
    .io_ho_out(bc_pe_197_io_ho_out),
    .io_res_out(bc_pe_197_io_res_out)
  );
  bc_pe bc_pe_198 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_198_clock),
    .reset(bc_pe_198_reset),
    .io_ho_input(bc_pe_198_io_ho_input),
    .io_ve_input(bc_pe_198_io_ve_input),
    .io_input_valid(bc_pe_198_io_input_valid),
    .io_iormac(bc_pe_198_io_iormac),
    .io_ve_out(bc_pe_198_io_ve_out),
    .io_ho_out(bc_pe_198_io_ho_out),
    .io_res_out(bc_pe_198_io_res_out)
  );
  bc_pe bc_pe_199 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_199_clock),
    .reset(bc_pe_199_reset),
    .io_ho_input(bc_pe_199_io_ho_input),
    .io_ve_input(bc_pe_199_io_ve_input),
    .io_input_valid(bc_pe_199_io_input_valid),
    .io_iormac(bc_pe_199_io_iormac),
    .io_ve_out(bc_pe_199_io_ve_out),
    .io_ho_out(bc_pe_199_io_ho_out),
    .io_res_out(bc_pe_199_io_res_out)
  );
  bc_pe bc_pe_200 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_200_clock),
    .reset(bc_pe_200_reset),
    .io_ho_input(bc_pe_200_io_ho_input),
    .io_ve_input(bc_pe_200_io_ve_input),
    .io_input_valid(bc_pe_200_io_input_valid),
    .io_iormac(bc_pe_200_io_iormac),
    .io_ve_out(bc_pe_200_io_ve_out),
    .io_ho_out(bc_pe_200_io_ho_out),
    .io_res_out(bc_pe_200_io_res_out)
  );
  bc_pe bc_pe_201 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_201_clock),
    .reset(bc_pe_201_reset),
    .io_ho_input(bc_pe_201_io_ho_input),
    .io_ve_input(bc_pe_201_io_ve_input),
    .io_input_valid(bc_pe_201_io_input_valid),
    .io_iormac(bc_pe_201_io_iormac),
    .io_ve_out(bc_pe_201_io_ve_out),
    .io_ho_out(bc_pe_201_io_ho_out),
    .io_res_out(bc_pe_201_io_res_out)
  );
  bc_pe bc_pe_202 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_202_clock),
    .reset(bc_pe_202_reset),
    .io_ho_input(bc_pe_202_io_ho_input),
    .io_ve_input(bc_pe_202_io_ve_input),
    .io_input_valid(bc_pe_202_io_input_valid),
    .io_iormac(bc_pe_202_io_iormac),
    .io_ve_out(bc_pe_202_io_ve_out),
    .io_ho_out(bc_pe_202_io_ho_out),
    .io_res_out(bc_pe_202_io_res_out)
  );
  bc_pe bc_pe_203 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_203_clock),
    .reset(bc_pe_203_reset),
    .io_ho_input(bc_pe_203_io_ho_input),
    .io_ve_input(bc_pe_203_io_ve_input),
    .io_input_valid(bc_pe_203_io_input_valid),
    .io_iormac(bc_pe_203_io_iormac),
    .io_ve_out(bc_pe_203_io_ve_out),
    .io_ho_out(bc_pe_203_io_ho_out),
    .io_res_out(bc_pe_203_io_res_out)
  );
  bc_pe bc_pe_204 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_204_clock),
    .reset(bc_pe_204_reset),
    .io_ho_input(bc_pe_204_io_ho_input),
    .io_ve_input(bc_pe_204_io_ve_input),
    .io_input_valid(bc_pe_204_io_input_valid),
    .io_iormac(bc_pe_204_io_iormac),
    .io_ve_out(bc_pe_204_io_ve_out),
    .io_ho_out(bc_pe_204_io_ho_out),
    .io_res_out(bc_pe_204_io_res_out)
  );
  bc_pe bc_pe_205 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_205_clock),
    .reset(bc_pe_205_reset),
    .io_ho_input(bc_pe_205_io_ho_input),
    .io_ve_input(bc_pe_205_io_ve_input),
    .io_input_valid(bc_pe_205_io_input_valid),
    .io_iormac(bc_pe_205_io_iormac),
    .io_ve_out(bc_pe_205_io_ve_out),
    .io_ho_out(bc_pe_205_io_ho_out),
    .io_res_out(bc_pe_205_io_res_out)
  );
  bc_pe bc_pe_206 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_206_clock),
    .reset(bc_pe_206_reset),
    .io_ho_input(bc_pe_206_io_ho_input),
    .io_ve_input(bc_pe_206_io_ve_input),
    .io_input_valid(bc_pe_206_io_input_valid),
    .io_iormac(bc_pe_206_io_iormac),
    .io_ve_out(bc_pe_206_io_ve_out),
    .io_ho_out(bc_pe_206_io_ho_out),
    .io_res_out(bc_pe_206_io_res_out)
  );
  bc_pe bc_pe_207 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_207_clock),
    .reset(bc_pe_207_reset),
    .io_ho_input(bc_pe_207_io_ho_input),
    .io_ve_input(bc_pe_207_io_ve_input),
    .io_input_valid(bc_pe_207_io_input_valid),
    .io_iormac(bc_pe_207_io_iormac),
    .io_ve_out(bc_pe_207_io_ve_out),
    .io_ho_out(bc_pe_207_io_ho_out),
    .io_res_out(bc_pe_207_io_res_out)
  );
  bc_pe bc_pe_208 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_208_clock),
    .reset(bc_pe_208_reset),
    .io_ho_input(bc_pe_208_io_ho_input),
    .io_ve_input(bc_pe_208_io_ve_input),
    .io_input_valid(bc_pe_208_io_input_valid),
    .io_iormac(bc_pe_208_io_iormac),
    .io_ve_out(bc_pe_208_io_ve_out),
    .io_ho_out(bc_pe_208_io_ho_out),
    .io_res_out(bc_pe_208_io_res_out)
  );
  bc_pe bc_pe_209 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_209_clock),
    .reset(bc_pe_209_reset),
    .io_ho_input(bc_pe_209_io_ho_input),
    .io_ve_input(bc_pe_209_io_ve_input),
    .io_input_valid(bc_pe_209_io_input_valid),
    .io_iormac(bc_pe_209_io_iormac),
    .io_ve_out(bc_pe_209_io_ve_out),
    .io_ho_out(bc_pe_209_io_ho_out),
    .io_res_out(bc_pe_209_io_res_out)
  );
  bc_pe bc_pe_210 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_210_clock),
    .reset(bc_pe_210_reset),
    .io_ho_input(bc_pe_210_io_ho_input),
    .io_ve_input(bc_pe_210_io_ve_input),
    .io_input_valid(bc_pe_210_io_input_valid),
    .io_iormac(bc_pe_210_io_iormac),
    .io_ve_out(bc_pe_210_io_ve_out),
    .io_ho_out(bc_pe_210_io_ho_out),
    .io_res_out(bc_pe_210_io_res_out)
  );
  bc_pe bc_pe_211 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_211_clock),
    .reset(bc_pe_211_reset),
    .io_ho_input(bc_pe_211_io_ho_input),
    .io_ve_input(bc_pe_211_io_ve_input),
    .io_input_valid(bc_pe_211_io_input_valid),
    .io_iormac(bc_pe_211_io_iormac),
    .io_ve_out(bc_pe_211_io_ve_out),
    .io_ho_out(bc_pe_211_io_ho_out),
    .io_res_out(bc_pe_211_io_res_out)
  );
  bc_pe bc_pe_212 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_212_clock),
    .reset(bc_pe_212_reset),
    .io_ho_input(bc_pe_212_io_ho_input),
    .io_ve_input(bc_pe_212_io_ve_input),
    .io_input_valid(bc_pe_212_io_input_valid),
    .io_iormac(bc_pe_212_io_iormac),
    .io_ve_out(bc_pe_212_io_ve_out),
    .io_ho_out(bc_pe_212_io_ho_out),
    .io_res_out(bc_pe_212_io_res_out)
  );
  bc_pe bc_pe_213 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_213_clock),
    .reset(bc_pe_213_reset),
    .io_ho_input(bc_pe_213_io_ho_input),
    .io_ve_input(bc_pe_213_io_ve_input),
    .io_input_valid(bc_pe_213_io_input_valid),
    .io_iormac(bc_pe_213_io_iormac),
    .io_ve_out(bc_pe_213_io_ve_out),
    .io_ho_out(bc_pe_213_io_ho_out),
    .io_res_out(bc_pe_213_io_res_out)
  );
  bc_pe bc_pe_214 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_214_clock),
    .reset(bc_pe_214_reset),
    .io_ho_input(bc_pe_214_io_ho_input),
    .io_ve_input(bc_pe_214_io_ve_input),
    .io_input_valid(bc_pe_214_io_input_valid),
    .io_iormac(bc_pe_214_io_iormac),
    .io_ve_out(bc_pe_214_io_ve_out),
    .io_ho_out(bc_pe_214_io_ho_out),
    .io_res_out(bc_pe_214_io_res_out)
  );
  bc_pe bc_pe_215 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_215_clock),
    .reset(bc_pe_215_reset),
    .io_ho_input(bc_pe_215_io_ho_input),
    .io_ve_input(bc_pe_215_io_ve_input),
    .io_input_valid(bc_pe_215_io_input_valid),
    .io_iormac(bc_pe_215_io_iormac),
    .io_ve_out(bc_pe_215_io_ve_out),
    .io_ho_out(bc_pe_215_io_ho_out),
    .io_res_out(bc_pe_215_io_res_out)
  );
  bc_pe bc_pe_216 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_216_clock),
    .reset(bc_pe_216_reset),
    .io_ho_input(bc_pe_216_io_ho_input),
    .io_ve_input(bc_pe_216_io_ve_input),
    .io_input_valid(bc_pe_216_io_input_valid),
    .io_iormac(bc_pe_216_io_iormac),
    .io_ve_out(bc_pe_216_io_ve_out),
    .io_ho_out(bc_pe_216_io_ho_out),
    .io_res_out(bc_pe_216_io_res_out)
  );
  bc_pe bc_pe_217 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_217_clock),
    .reset(bc_pe_217_reset),
    .io_ho_input(bc_pe_217_io_ho_input),
    .io_ve_input(bc_pe_217_io_ve_input),
    .io_input_valid(bc_pe_217_io_input_valid),
    .io_iormac(bc_pe_217_io_iormac),
    .io_ve_out(bc_pe_217_io_ve_out),
    .io_ho_out(bc_pe_217_io_ho_out),
    .io_res_out(bc_pe_217_io_res_out)
  );
  bc_pe bc_pe_218 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_218_clock),
    .reset(bc_pe_218_reset),
    .io_ho_input(bc_pe_218_io_ho_input),
    .io_ve_input(bc_pe_218_io_ve_input),
    .io_input_valid(bc_pe_218_io_input_valid),
    .io_iormac(bc_pe_218_io_iormac),
    .io_ve_out(bc_pe_218_io_ve_out),
    .io_ho_out(bc_pe_218_io_ho_out),
    .io_res_out(bc_pe_218_io_res_out)
  );
  bc_pe bc_pe_219 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_219_clock),
    .reset(bc_pe_219_reset),
    .io_ho_input(bc_pe_219_io_ho_input),
    .io_ve_input(bc_pe_219_io_ve_input),
    .io_input_valid(bc_pe_219_io_input_valid),
    .io_iormac(bc_pe_219_io_iormac),
    .io_ve_out(bc_pe_219_io_ve_out),
    .io_ho_out(bc_pe_219_io_ho_out),
    .io_res_out(bc_pe_219_io_res_out)
  );
  bc_pe bc_pe_220 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_220_clock),
    .reset(bc_pe_220_reset),
    .io_ho_input(bc_pe_220_io_ho_input),
    .io_ve_input(bc_pe_220_io_ve_input),
    .io_input_valid(bc_pe_220_io_input_valid),
    .io_iormac(bc_pe_220_io_iormac),
    .io_ve_out(bc_pe_220_io_ve_out),
    .io_ho_out(bc_pe_220_io_ho_out),
    .io_res_out(bc_pe_220_io_res_out)
  );
  bc_pe bc_pe_221 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_221_clock),
    .reset(bc_pe_221_reset),
    .io_ho_input(bc_pe_221_io_ho_input),
    .io_ve_input(bc_pe_221_io_ve_input),
    .io_input_valid(bc_pe_221_io_input_valid),
    .io_iormac(bc_pe_221_io_iormac),
    .io_ve_out(bc_pe_221_io_ve_out),
    .io_ho_out(bc_pe_221_io_ho_out),
    .io_res_out(bc_pe_221_io_res_out)
  );
  bc_pe bc_pe_222 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_222_clock),
    .reset(bc_pe_222_reset),
    .io_ho_input(bc_pe_222_io_ho_input),
    .io_ve_input(bc_pe_222_io_ve_input),
    .io_input_valid(bc_pe_222_io_input_valid),
    .io_iormac(bc_pe_222_io_iormac),
    .io_ve_out(bc_pe_222_io_ve_out),
    .io_ho_out(bc_pe_222_io_ho_out),
    .io_res_out(bc_pe_222_io_res_out)
  );
  bc_pe bc_pe_223 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_223_clock),
    .reset(bc_pe_223_reset),
    .io_ho_input(bc_pe_223_io_ho_input),
    .io_ve_input(bc_pe_223_io_ve_input),
    .io_input_valid(bc_pe_223_io_input_valid),
    .io_iormac(bc_pe_223_io_iormac),
    .io_ve_out(bc_pe_223_io_ve_out),
    .io_ho_out(bc_pe_223_io_ho_out),
    .io_res_out(bc_pe_223_io_res_out)
  );
  bc_pe bc_pe_224 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_224_clock),
    .reset(bc_pe_224_reset),
    .io_ho_input(bc_pe_224_io_ho_input),
    .io_ve_input(bc_pe_224_io_ve_input),
    .io_input_valid(bc_pe_224_io_input_valid),
    .io_iormac(bc_pe_224_io_iormac),
    .io_ve_out(bc_pe_224_io_ve_out),
    .io_ho_out(bc_pe_224_io_ho_out),
    .io_res_out(bc_pe_224_io_res_out)
  );
  bc_pe bc_pe_225 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_225_clock),
    .reset(bc_pe_225_reset),
    .io_ho_input(bc_pe_225_io_ho_input),
    .io_ve_input(bc_pe_225_io_ve_input),
    .io_input_valid(bc_pe_225_io_input_valid),
    .io_iormac(bc_pe_225_io_iormac),
    .io_ve_out(bc_pe_225_io_ve_out),
    .io_ho_out(bc_pe_225_io_ho_out),
    .io_res_out(bc_pe_225_io_res_out)
  );
  bc_pe bc_pe_226 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_226_clock),
    .reset(bc_pe_226_reset),
    .io_ho_input(bc_pe_226_io_ho_input),
    .io_ve_input(bc_pe_226_io_ve_input),
    .io_input_valid(bc_pe_226_io_input_valid),
    .io_iormac(bc_pe_226_io_iormac),
    .io_ve_out(bc_pe_226_io_ve_out),
    .io_ho_out(bc_pe_226_io_ho_out),
    .io_res_out(bc_pe_226_io_res_out)
  );
  bc_pe bc_pe_227 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_227_clock),
    .reset(bc_pe_227_reset),
    .io_ho_input(bc_pe_227_io_ho_input),
    .io_ve_input(bc_pe_227_io_ve_input),
    .io_input_valid(bc_pe_227_io_input_valid),
    .io_iormac(bc_pe_227_io_iormac),
    .io_ve_out(bc_pe_227_io_ve_out),
    .io_ho_out(bc_pe_227_io_ho_out),
    .io_res_out(bc_pe_227_io_res_out)
  );
  bc_pe bc_pe_228 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_228_clock),
    .reset(bc_pe_228_reset),
    .io_ho_input(bc_pe_228_io_ho_input),
    .io_ve_input(bc_pe_228_io_ve_input),
    .io_input_valid(bc_pe_228_io_input_valid),
    .io_iormac(bc_pe_228_io_iormac),
    .io_ve_out(bc_pe_228_io_ve_out),
    .io_ho_out(bc_pe_228_io_ho_out),
    .io_res_out(bc_pe_228_io_res_out)
  );
  bc_pe bc_pe_229 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_229_clock),
    .reset(bc_pe_229_reset),
    .io_ho_input(bc_pe_229_io_ho_input),
    .io_ve_input(bc_pe_229_io_ve_input),
    .io_input_valid(bc_pe_229_io_input_valid),
    .io_iormac(bc_pe_229_io_iormac),
    .io_ve_out(bc_pe_229_io_ve_out),
    .io_ho_out(bc_pe_229_io_ho_out),
    .io_res_out(bc_pe_229_io_res_out)
  );
  bc_pe bc_pe_230 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_230_clock),
    .reset(bc_pe_230_reset),
    .io_ho_input(bc_pe_230_io_ho_input),
    .io_ve_input(bc_pe_230_io_ve_input),
    .io_input_valid(bc_pe_230_io_input_valid),
    .io_iormac(bc_pe_230_io_iormac),
    .io_ve_out(bc_pe_230_io_ve_out),
    .io_ho_out(bc_pe_230_io_ho_out),
    .io_res_out(bc_pe_230_io_res_out)
  );
  bc_pe bc_pe_231 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_231_clock),
    .reset(bc_pe_231_reset),
    .io_ho_input(bc_pe_231_io_ho_input),
    .io_ve_input(bc_pe_231_io_ve_input),
    .io_input_valid(bc_pe_231_io_input_valid),
    .io_iormac(bc_pe_231_io_iormac),
    .io_ve_out(bc_pe_231_io_ve_out),
    .io_ho_out(bc_pe_231_io_ho_out),
    .io_res_out(bc_pe_231_io_res_out)
  );
  bc_pe bc_pe_232 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_232_clock),
    .reset(bc_pe_232_reset),
    .io_ho_input(bc_pe_232_io_ho_input),
    .io_ve_input(bc_pe_232_io_ve_input),
    .io_input_valid(bc_pe_232_io_input_valid),
    .io_iormac(bc_pe_232_io_iormac),
    .io_ve_out(bc_pe_232_io_ve_out),
    .io_ho_out(bc_pe_232_io_ho_out),
    .io_res_out(bc_pe_232_io_res_out)
  );
  bc_pe bc_pe_233 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_233_clock),
    .reset(bc_pe_233_reset),
    .io_ho_input(bc_pe_233_io_ho_input),
    .io_ve_input(bc_pe_233_io_ve_input),
    .io_input_valid(bc_pe_233_io_input_valid),
    .io_iormac(bc_pe_233_io_iormac),
    .io_ve_out(bc_pe_233_io_ve_out),
    .io_ho_out(bc_pe_233_io_ho_out),
    .io_res_out(bc_pe_233_io_res_out)
  );
  bc_pe bc_pe_234 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_234_clock),
    .reset(bc_pe_234_reset),
    .io_ho_input(bc_pe_234_io_ho_input),
    .io_ve_input(bc_pe_234_io_ve_input),
    .io_input_valid(bc_pe_234_io_input_valid),
    .io_iormac(bc_pe_234_io_iormac),
    .io_ve_out(bc_pe_234_io_ve_out),
    .io_ho_out(bc_pe_234_io_ho_out),
    .io_res_out(bc_pe_234_io_res_out)
  );
  bc_pe bc_pe_235 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_235_clock),
    .reset(bc_pe_235_reset),
    .io_ho_input(bc_pe_235_io_ho_input),
    .io_ve_input(bc_pe_235_io_ve_input),
    .io_input_valid(bc_pe_235_io_input_valid),
    .io_iormac(bc_pe_235_io_iormac),
    .io_ve_out(bc_pe_235_io_ve_out),
    .io_ho_out(bc_pe_235_io_ho_out),
    .io_res_out(bc_pe_235_io_res_out)
  );
  bc_pe bc_pe_236 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_236_clock),
    .reset(bc_pe_236_reset),
    .io_ho_input(bc_pe_236_io_ho_input),
    .io_ve_input(bc_pe_236_io_ve_input),
    .io_input_valid(bc_pe_236_io_input_valid),
    .io_iormac(bc_pe_236_io_iormac),
    .io_ve_out(bc_pe_236_io_ve_out),
    .io_ho_out(bc_pe_236_io_ho_out),
    .io_res_out(bc_pe_236_io_res_out)
  );
  bc_pe bc_pe_237 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_237_clock),
    .reset(bc_pe_237_reset),
    .io_ho_input(bc_pe_237_io_ho_input),
    .io_ve_input(bc_pe_237_io_ve_input),
    .io_input_valid(bc_pe_237_io_input_valid),
    .io_iormac(bc_pe_237_io_iormac),
    .io_ve_out(bc_pe_237_io_ve_out),
    .io_ho_out(bc_pe_237_io_ho_out),
    .io_res_out(bc_pe_237_io_res_out)
  );
  bc_pe bc_pe_238 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_238_clock),
    .reset(bc_pe_238_reset),
    .io_ho_input(bc_pe_238_io_ho_input),
    .io_ve_input(bc_pe_238_io_ve_input),
    .io_input_valid(bc_pe_238_io_input_valid),
    .io_iormac(bc_pe_238_io_iormac),
    .io_ve_out(bc_pe_238_io_ve_out),
    .io_ho_out(bc_pe_238_io_ho_out),
    .io_res_out(bc_pe_238_io_res_out)
  );
  bc_pe bc_pe_239 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_239_clock),
    .reset(bc_pe_239_reset),
    .io_ho_input(bc_pe_239_io_ho_input),
    .io_ve_input(bc_pe_239_io_ve_input),
    .io_input_valid(bc_pe_239_io_input_valid),
    .io_iormac(bc_pe_239_io_iormac),
    .io_ve_out(bc_pe_239_io_ve_out),
    .io_ho_out(bc_pe_239_io_ho_out),
    .io_res_out(bc_pe_239_io_res_out)
  );
  bc_pe bc_pe_240 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_240_clock),
    .reset(bc_pe_240_reset),
    .io_ho_input(bc_pe_240_io_ho_input),
    .io_ve_input(bc_pe_240_io_ve_input),
    .io_input_valid(bc_pe_240_io_input_valid),
    .io_iormac(bc_pe_240_io_iormac),
    .io_ve_out(bc_pe_240_io_ve_out),
    .io_ho_out(bc_pe_240_io_ho_out),
    .io_res_out(bc_pe_240_io_res_out)
  );
  bc_pe bc_pe_241 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_241_clock),
    .reset(bc_pe_241_reset),
    .io_ho_input(bc_pe_241_io_ho_input),
    .io_ve_input(bc_pe_241_io_ve_input),
    .io_input_valid(bc_pe_241_io_input_valid),
    .io_iormac(bc_pe_241_io_iormac),
    .io_ve_out(bc_pe_241_io_ve_out),
    .io_ho_out(bc_pe_241_io_ho_out),
    .io_res_out(bc_pe_241_io_res_out)
  );
  bc_pe bc_pe_242 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_242_clock),
    .reset(bc_pe_242_reset),
    .io_ho_input(bc_pe_242_io_ho_input),
    .io_ve_input(bc_pe_242_io_ve_input),
    .io_input_valid(bc_pe_242_io_input_valid),
    .io_iormac(bc_pe_242_io_iormac),
    .io_ve_out(bc_pe_242_io_ve_out),
    .io_ho_out(bc_pe_242_io_ho_out),
    .io_res_out(bc_pe_242_io_res_out)
  );
  bc_pe bc_pe_243 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_243_clock),
    .reset(bc_pe_243_reset),
    .io_ho_input(bc_pe_243_io_ho_input),
    .io_ve_input(bc_pe_243_io_ve_input),
    .io_input_valid(bc_pe_243_io_input_valid),
    .io_iormac(bc_pe_243_io_iormac),
    .io_ve_out(bc_pe_243_io_ve_out),
    .io_ho_out(bc_pe_243_io_ho_out),
    .io_res_out(bc_pe_243_io_res_out)
  );
  bc_pe bc_pe_244 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_244_clock),
    .reset(bc_pe_244_reset),
    .io_ho_input(bc_pe_244_io_ho_input),
    .io_ve_input(bc_pe_244_io_ve_input),
    .io_input_valid(bc_pe_244_io_input_valid),
    .io_iormac(bc_pe_244_io_iormac),
    .io_ve_out(bc_pe_244_io_ve_out),
    .io_ho_out(bc_pe_244_io_ho_out),
    .io_res_out(bc_pe_244_io_res_out)
  );
  bc_pe bc_pe_245 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_245_clock),
    .reset(bc_pe_245_reset),
    .io_ho_input(bc_pe_245_io_ho_input),
    .io_ve_input(bc_pe_245_io_ve_input),
    .io_input_valid(bc_pe_245_io_input_valid),
    .io_iormac(bc_pe_245_io_iormac),
    .io_ve_out(bc_pe_245_io_ve_out),
    .io_ho_out(bc_pe_245_io_ho_out),
    .io_res_out(bc_pe_245_io_res_out)
  );
  bc_pe bc_pe_246 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_246_clock),
    .reset(bc_pe_246_reset),
    .io_ho_input(bc_pe_246_io_ho_input),
    .io_ve_input(bc_pe_246_io_ve_input),
    .io_input_valid(bc_pe_246_io_input_valid),
    .io_iormac(bc_pe_246_io_iormac),
    .io_ve_out(bc_pe_246_io_ve_out),
    .io_ho_out(bc_pe_246_io_ho_out),
    .io_res_out(bc_pe_246_io_res_out)
  );
  bc_pe bc_pe_247 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_247_clock),
    .reset(bc_pe_247_reset),
    .io_ho_input(bc_pe_247_io_ho_input),
    .io_ve_input(bc_pe_247_io_ve_input),
    .io_input_valid(bc_pe_247_io_input_valid),
    .io_iormac(bc_pe_247_io_iormac),
    .io_ve_out(bc_pe_247_io_ve_out),
    .io_ho_out(bc_pe_247_io_ho_out),
    .io_res_out(bc_pe_247_io_res_out)
  );
  bc_pe bc_pe_248 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_248_clock),
    .reset(bc_pe_248_reset),
    .io_ho_input(bc_pe_248_io_ho_input),
    .io_ve_input(bc_pe_248_io_ve_input),
    .io_input_valid(bc_pe_248_io_input_valid),
    .io_iormac(bc_pe_248_io_iormac),
    .io_ve_out(bc_pe_248_io_ve_out),
    .io_ho_out(bc_pe_248_io_ho_out),
    .io_res_out(bc_pe_248_io_res_out)
  );
  bc_pe bc_pe_249 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_249_clock),
    .reset(bc_pe_249_reset),
    .io_ho_input(bc_pe_249_io_ho_input),
    .io_ve_input(bc_pe_249_io_ve_input),
    .io_input_valid(bc_pe_249_io_input_valid),
    .io_iormac(bc_pe_249_io_iormac),
    .io_ve_out(bc_pe_249_io_ve_out),
    .io_ho_out(bc_pe_249_io_ho_out),
    .io_res_out(bc_pe_249_io_res_out)
  );
  bc_pe bc_pe_250 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_250_clock),
    .reset(bc_pe_250_reset),
    .io_ho_input(bc_pe_250_io_ho_input),
    .io_ve_input(bc_pe_250_io_ve_input),
    .io_input_valid(bc_pe_250_io_input_valid),
    .io_iormac(bc_pe_250_io_iormac),
    .io_ve_out(bc_pe_250_io_ve_out),
    .io_ho_out(bc_pe_250_io_ho_out),
    .io_res_out(bc_pe_250_io_res_out)
  );
  bc_pe bc_pe_251 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_251_clock),
    .reset(bc_pe_251_reset),
    .io_ho_input(bc_pe_251_io_ho_input),
    .io_ve_input(bc_pe_251_io_ve_input),
    .io_input_valid(bc_pe_251_io_input_valid),
    .io_iormac(bc_pe_251_io_iormac),
    .io_ve_out(bc_pe_251_io_ve_out),
    .io_ho_out(bc_pe_251_io_ho_out),
    .io_res_out(bc_pe_251_io_res_out)
  );
  bc_pe bc_pe_252 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_252_clock),
    .reset(bc_pe_252_reset),
    .io_ho_input(bc_pe_252_io_ho_input),
    .io_ve_input(bc_pe_252_io_ve_input),
    .io_input_valid(bc_pe_252_io_input_valid),
    .io_iormac(bc_pe_252_io_iormac),
    .io_ve_out(bc_pe_252_io_ve_out),
    .io_ho_out(bc_pe_252_io_ho_out),
    .io_res_out(bc_pe_252_io_res_out)
  );
  bc_pe bc_pe_253 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_253_clock),
    .reset(bc_pe_253_reset),
    .io_ho_input(bc_pe_253_io_ho_input),
    .io_ve_input(bc_pe_253_io_ve_input),
    .io_input_valid(bc_pe_253_io_input_valid),
    .io_iormac(bc_pe_253_io_iormac),
    .io_ve_out(bc_pe_253_io_ve_out),
    .io_ho_out(bc_pe_253_io_ho_out),
    .io_res_out(bc_pe_253_io_res_out)
  );
  bc_pe bc_pe_254 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_254_clock),
    .reset(bc_pe_254_reset),
    .io_ho_input(bc_pe_254_io_ho_input),
    .io_ve_input(bc_pe_254_io_ve_input),
    .io_input_valid(bc_pe_254_io_input_valid),
    .io_iormac(bc_pe_254_io_iormac),
    .io_ve_out(bc_pe_254_io_ve_out),
    .io_ho_out(bc_pe_254_io_ho_out),
    .io_res_out(bc_pe_254_io_res_out)
  );
  bc_pe bc_pe_255 ( // @[bc_mmul.scala 23:11]
    .clock(bc_pe_255_clock),
    .reset(bc_pe_255_reset),
    .io_ho_input(bc_pe_255_io_ho_input),
    .io_ve_input(bc_pe_255_io_ve_input),
    .io_input_valid(bc_pe_255_io_input_valid),
    .io_iormac(bc_pe_255_io_iormac),
    .io_ve_out(bc_pe_255_io_ve_out),
    .io_ho_out(bc_pe_255_io_ho_out),
    .io_res_out(bc_pe_255_io_res_out)
  );
  assign io_out_0 = bc_pe_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_1 = bc_pe_1_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_2 = bc_pe_2_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_3 = bc_pe_3_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_4 = bc_pe_4_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_5 = bc_pe_5_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_6 = bc_pe_6_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_7 = bc_pe_7_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_8 = bc_pe_8_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_9 = bc_pe_9_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_10 = bc_pe_10_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_11 = bc_pe_11_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_12 = bc_pe_12_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_13 = bc_pe_13_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_14 = bc_pe_14_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_15 = bc_pe_15_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_16 = bc_pe_16_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_17 = bc_pe_17_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_18 = bc_pe_18_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_19 = bc_pe_19_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_20 = bc_pe_20_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_21 = bc_pe_21_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_22 = bc_pe_22_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_23 = bc_pe_23_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_24 = bc_pe_24_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_25 = bc_pe_25_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_26 = bc_pe_26_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_27 = bc_pe_27_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_28 = bc_pe_28_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_29 = bc_pe_29_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_30 = bc_pe_30_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_31 = bc_pe_31_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_32 = bc_pe_32_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_33 = bc_pe_33_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_34 = bc_pe_34_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_35 = bc_pe_35_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_36 = bc_pe_36_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_37 = bc_pe_37_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_38 = bc_pe_38_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_39 = bc_pe_39_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_40 = bc_pe_40_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_41 = bc_pe_41_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_42 = bc_pe_42_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_43 = bc_pe_43_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_44 = bc_pe_44_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_45 = bc_pe_45_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_46 = bc_pe_46_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_47 = bc_pe_47_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_48 = bc_pe_48_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_49 = bc_pe_49_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_50 = bc_pe_50_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_51 = bc_pe_51_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_52 = bc_pe_52_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_53 = bc_pe_53_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_54 = bc_pe_54_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_55 = bc_pe_55_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_56 = bc_pe_56_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_57 = bc_pe_57_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_58 = bc_pe_58_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_59 = bc_pe_59_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_60 = bc_pe_60_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_61 = bc_pe_61_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_62 = bc_pe_62_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_63 = bc_pe_63_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_64 = bc_pe_64_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_65 = bc_pe_65_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_66 = bc_pe_66_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_67 = bc_pe_67_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_68 = bc_pe_68_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_69 = bc_pe_69_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_70 = bc_pe_70_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_71 = bc_pe_71_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_72 = bc_pe_72_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_73 = bc_pe_73_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_74 = bc_pe_74_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_75 = bc_pe_75_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_76 = bc_pe_76_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_77 = bc_pe_77_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_78 = bc_pe_78_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_79 = bc_pe_79_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_80 = bc_pe_80_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_81 = bc_pe_81_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_82 = bc_pe_82_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_83 = bc_pe_83_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_84 = bc_pe_84_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_85 = bc_pe_85_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_86 = bc_pe_86_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_87 = bc_pe_87_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_88 = bc_pe_88_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_89 = bc_pe_89_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_90 = bc_pe_90_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_91 = bc_pe_91_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_92 = bc_pe_92_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_93 = bc_pe_93_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_94 = bc_pe_94_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_95 = bc_pe_95_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_96 = bc_pe_96_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_97 = bc_pe_97_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_98 = bc_pe_98_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_99 = bc_pe_99_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_100 = bc_pe_100_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_101 = bc_pe_101_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_102 = bc_pe_102_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_103 = bc_pe_103_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_104 = bc_pe_104_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_105 = bc_pe_105_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_106 = bc_pe_106_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_107 = bc_pe_107_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_108 = bc_pe_108_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_109 = bc_pe_109_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_110 = bc_pe_110_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_111 = bc_pe_111_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_112 = bc_pe_112_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_113 = bc_pe_113_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_114 = bc_pe_114_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_115 = bc_pe_115_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_116 = bc_pe_116_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_117 = bc_pe_117_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_118 = bc_pe_118_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_119 = bc_pe_119_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_120 = bc_pe_120_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_121 = bc_pe_121_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_122 = bc_pe_122_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_123 = bc_pe_123_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_124 = bc_pe_124_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_125 = bc_pe_125_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_126 = bc_pe_126_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_127 = bc_pe_127_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_128 = bc_pe_128_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_129 = bc_pe_129_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_130 = bc_pe_130_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_131 = bc_pe_131_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_132 = bc_pe_132_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_133 = bc_pe_133_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_134 = bc_pe_134_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_135 = bc_pe_135_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_136 = bc_pe_136_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_137 = bc_pe_137_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_138 = bc_pe_138_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_139 = bc_pe_139_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_140 = bc_pe_140_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_141 = bc_pe_141_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_142 = bc_pe_142_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_143 = bc_pe_143_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_144 = bc_pe_144_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_145 = bc_pe_145_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_146 = bc_pe_146_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_147 = bc_pe_147_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_148 = bc_pe_148_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_149 = bc_pe_149_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_150 = bc_pe_150_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_151 = bc_pe_151_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_152 = bc_pe_152_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_153 = bc_pe_153_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_154 = bc_pe_154_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_155 = bc_pe_155_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_156 = bc_pe_156_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_157 = bc_pe_157_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_158 = bc_pe_158_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_159 = bc_pe_159_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_160 = bc_pe_160_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_161 = bc_pe_161_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_162 = bc_pe_162_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_163 = bc_pe_163_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_164 = bc_pe_164_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_165 = bc_pe_165_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_166 = bc_pe_166_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_167 = bc_pe_167_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_168 = bc_pe_168_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_169 = bc_pe_169_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_170 = bc_pe_170_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_171 = bc_pe_171_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_172 = bc_pe_172_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_173 = bc_pe_173_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_174 = bc_pe_174_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_175 = bc_pe_175_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_176 = bc_pe_176_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_177 = bc_pe_177_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_178 = bc_pe_178_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_179 = bc_pe_179_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_180 = bc_pe_180_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_181 = bc_pe_181_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_182 = bc_pe_182_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_183 = bc_pe_183_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_184 = bc_pe_184_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_185 = bc_pe_185_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_186 = bc_pe_186_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_187 = bc_pe_187_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_188 = bc_pe_188_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_189 = bc_pe_189_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_190 = bc_pe_190_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_191 = bc_pe_191_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_192 = bc_pe_192_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_193 = bc_pe_193_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_194 = bc_pe_194_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_195 = bc_pe_195_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_196 = bc_pe_196_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_197 = bc_pe_197_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_198 = bc_pe_198_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_199 = bc_pe_199_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_200 = bc_pe_200_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_201 = bc_pe_201_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_202 = bc_pe_202_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_203 = bc_pe_203_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_204 = bc_pe_204_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_205 = bc_pe_205_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_206 = bc_pe_206_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_207 = bc_pe_207_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_208 = bc_pe_208_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_209 = bc_pe_209_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_210 = bc_pe_210_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_211 = bc_pe_211_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_212 = bc_pe_212_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_213 = bc_pe_213_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_214 = bc_pe_214_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_215 = bc_pe_215_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_216 = bc_pe_216_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_217 = bc_pe_217_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_218 = bc_pe_218_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_219 = bc_pe_219_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_220 = bc_pe_220_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_221 = bc_pe_221_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_222 = bc_pe_222_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_223 = bc_pe_223_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_224 = bc_pe_224_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_225 = bc_pe_225_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_226 = bc_pe_226_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_227 = bc_pe_227_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_228 = bc_pe_228_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_229 = bc_pe_229_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_230 = bc_pe_230_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_231 = bc_pe_231_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_232 = bc_pe_232_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_233 = bc_pe_233_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_234 = bc_pe_234_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_235 = bc_pe_235_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_236 = bc_pe_236_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_237 = bc_pe_237_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_238 = bc_pe_238_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_239 = bc_pe_239_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_240 = bc_pe_240_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_241 = bc_pe_241_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_242 = bc_pe_242_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_243 = bc_pe_243_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_244 = bc_pe_244_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_245 = bc_pe_245_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_246 = bc_pe_246_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_247 = bc_pe_247_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_248 = bc_pe_248_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_249 = bc_pe_249_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_250 = bc_pe_250_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_251 = bc_pe_251_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_252 = bc_pe_252_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_253 = bc_pe_253_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_254 = bc_pe_254_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign io_out_255 = bc_pe_255_io_res_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_clock = clock;
  assign bc_pe_reset = reset;
  assign bc_pe_io_ho_input = io_x_input_0; // @[bc_mmul.scala 22:28 38:42]
  assign bc_pe_io_ve_input = io_w_input_0; // @[bc_mmul.scala 22:28 37:42]
  assign bc_pe_io_input_valid = io_input_valid_0; // @[bc_mmul.scala 22:28 39:42]
  assign bc_pe_io_iormac = io_iormac_0; // @[bc_mmul.scala 22:28 40:42]
  assign bc_pe_1_clock = clock;
  assign bc_pe_1_reset = reset;
  assign bc_pe_1_io_ho_input = bc_pe_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_1_io_ve_input = io_w_input_1; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_1_io_input_valid = io_input_valid_1; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_1_io_iormac = io_iormac_1; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_2_clock = clock;
  assign bc_pe_2_reset = reset;
  assign bc_pe_2_io_ho_input = bc_pe_1_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_2_io_ve_input = io_w_input_2; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_2_io_input_valid = io_input_valid_2; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_2_io_iormac = io_iormac_2; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_3_clock = clock;
  assign bc_pe_3_reset = reset;
  assign bc_pe_3_io_ho_input = bc_pe_2_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_3_io_ve_input = io_w_input_3; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_3_io_input_valid = io_input_valid_3; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_3_io_iormac = io_iormac_3; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_4_clock = clock;
  assign bc_pe_4_reset = reset;
  assign bc_pe_4_io_ho_input = bc_pe_3_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_4_io_ve_input = io_w_input_4; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_4_io_input_valid = io_input_valid_4; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_4_io_iormac = io_iormac_4; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_5_clock = clock;
  assign bc_pe_5_reset = reset;
  assign bc_pe_5_io_ho_input = bc_pe_4_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_5_io_ve_input = io_w_input_5; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_5_io_input_valid = io_input_valid_5; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_5_io_iormac = io_iormac_5; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_6_clock = clock;
  assign bc_pe_6_reset = reset;
  assign bc_pe_6_io_ho_input = bc_pe_5_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_6_io_ve_input = io_w_input_6; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_6_io_input_valid = io_input_valid_6; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_6_io_iormac = io_iormac_6; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_7_clock = clock;
  assign bc_pe_7_reset = reset;
  assign bc_pe_7_io_ho_input = bc_pe_6_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_7_io_ve_input = io_w_input_7; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_7_io_input_valid = io_input_valid_7; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_7_io_iormac = io_iormac_7; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_8_clock = clock;
  assign bc_pe_8_reset = reset;
  assign bc_pe_8_io_ho_input = bc_pe_7_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_8_io_ve_input = io_w_input_8; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_8_io_input_valid = io_input_valid_8; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_8_io_iormac = io_iormac_8; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_9_clock = clock;
  assign bc_pe_9_reset = reset;
  assign bc_pe_9_io_ho_input = bc_pe_8_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_9_io_ve_input = io_w_input_9; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_9_io_input_valid = io_input_valid_9; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_9_io_iormac = io_iormac_9; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_10_clock = clock;
  assign bc_pe_10_reset = reset;
  assign bc_pe_10_io_ho_input = bc_pe_9_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_10_io_ve_input = io_w_input_10; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_10_io_input_valid = io_input_valid_10; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_10_io_iormac = io_iormac_10; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_11_clock = clock;
  assign bc_pe_11_reset = reset;
  assign bc_pe_11_io_ho_input = bc_pe_10_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_11_io_ve_input = io_w_input_11; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_11_io_input_valid = io_input_valid_11; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_11_io_iormac = io_iormac_11; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_12_clock = clock;
  assign bc_pe_12_reset = reset;
  assign bc_pe_12_io_ho_input = bc_pe_11_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_12_io_ve_input = io_w_input_12; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_12_io_input_valid = io_input_valid_12; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_12_io_iormac = io_iormac_12; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_13_clock = clock;
  assign bc_pe_13_reset = reset;
  assign bc_pe_13_io_ho_input = bc_pe_12_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_13_io_ve_input = io_w_input_13; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_13_io_input_valid = io_input_valid_13; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_13_io_iormac = io_iormac_13; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_14_clock = clock;
  assign bc_pe_14_reset = reset;
  assign bc_pe_14_io_ho_input = bc_pe_13_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_14_io_ve_input = io_w_input_14; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_14_io_input_valid = io_input_valid_14; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_14_io_iormac = io_iormac_14; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_15_clock = clock;
  assign bc_pe_15_reset = reset;
  assign bc_pe_15_io_ho_input = bc_pe_14_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_15_io_ve_input = io_w_input_15; // @[bc_mmul.scala 22:28 48:43]
  assign bc_pe_15_io_input_valid = io_input_valid_15; // @[bc_mmul.scala 22:28 50:43]
  assign bc_pe_15_io_iormac = io_iormac_15; // @[bc_mmul.scala 22:28 51:43]
  assign bc_pe_16_clock = clock;
  assign bc_pe_16_reset = reset;
  assign bc_pe_16_io_ho_input = io_x_input_1; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_16_io_ve_input = bc_pe_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_16_io_input_valid = io_input_valid_16; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_16_io_iormac = io_iormac_16; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_17_clock = clock;
  assign bc_pe_17_reset = reset;
  assign bc_pe_17_io_ho_input = bc_pe_16_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_17_io_ve_input = bc_pe_1_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_17_io_input_valid = io_input_valid_17; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_17_io_iormac = io_iormac_17; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_18_clock = clock;
  assign bc_pe_18_reset = reset;
  assign bc_pe_18_io_ho_input = bc_pe_17_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_18_io_ve_input = bc_pe_2_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_18_io_input_valid = io_input_valid_18; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_18_io_iormac = io_iormac_18; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_19_clock = clock;
  assign bc_pe_19_reset = reset;
  assign bc_pe_19_io_ho_input = bc_pe_18_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_19_io_ve_input = bc_pe_3_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_19_io_input_valid = io_input_valid_19; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_19_io_iormac = io_iormac_19; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_20_clock = clock;
  assign bc_pe_20_reset = reset;
  assign bc_pe_20_io_ho_input = bc_pe_19_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_20_io_ve_input = bc_pe_4_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_20_io_input_valid = io_input_valid_20; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_20_io_iormac = io_iormac_20; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_21_clock = clock;
  assign bc_pe_21_reset = reset;
  assign bc_pe_21_io_ho_input = bc_pe_20_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_21_io_ve_input = bc_pe_5_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_21_io_input_valid = io_input_valid_21; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_21_io_iormac = io_iormac_21; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_22_clock = clock;
  assign bc_pe_22_reset = reset;
  assign bc_pe_22_io_ho_input = bc_pe_21_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_22_io_ve_input = bc_pe_6_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_22_io_input_valid = io_input_valid_22; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_22_io_iormac = io_iormac_22; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_23_clock = clock;
  assign bc_pe_23_reset = reset;
  assign bc_pe_23_io_ho_input = bc_pe_22_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_23_io_ve_input = bc_pe_7_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_23_io_input_valid = io_input_valid_23; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_23_io_iormac = io_iormac_23; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_24_clock = clock;
  assign bc_pe_24_reset = reset;
  assign bc_pe_24_io_ho_input = bc_pe_23_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_24_io_ve_input = bc_pe_8_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_24_io_input_valid = io_input_valid_24; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_24_io_iormac = io_iormac_24; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_25_clock = clock;
  assign bc_pe_25_reset = reset;
  assign bc_pe_25_io_ho_input = bc_pe_24_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_25_io_ve_input = bc_pe_9_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_25_io_input_valid = io_input_valid_25; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_25_io_iormac = io_iormac_25; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_26_clock = clock;
  assign bc_pe_26_reset = reset;
  assign bc_pe_26_io_ho_input = bc_pe_25_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_26_io_ve_input = bc_pe_10_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_26_io_input_valid = io_input_valid_26; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_26_io_iormac = io_iormac_26; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_27_clock = clock;
  assign bc_pe_27_reset = reset;
  assign bc_pe_27_io_ho_input = bc_pe_26_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_27_io_ve_input = bc_pe_11_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_27_io_input_valid = io_input_valid_27; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_27_io_iormac = io_iormac_27; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_28_clock = clock;
  assign bc_pe_28_reset = reset;
  assign bc_pe_28_io_ho_input = bc_pe_27_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_28_io_ve_input = bc_pe_12_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_28_io_input_valid = io_input_valid_28; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_28_io_iormac = io_iormac_28; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_29_clock = clock;
  assign bc_pe_29_reset = reset;
  assign bc_pe_29_io_ho_input = bc_pe_28_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_29_io_ve_input = bc_pe_13_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_29_io_input_valid = io_input_valid_29; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_29_io_iormac = io_iormac_29; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_30_clock = clock;
  assign bc_pe_30_reset = reset;
  assign bc_pe_30_io_ho_input = bc_pe_29_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_30_io_ve_input = bc_pe_14_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_30_io_input_valid = io_input_valid_30; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_30_io_iormac = io_iormac_30; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_31_clock = clock;
  assign bc_pe_31_reset = reset;
  assign bc_pe_31_io_ho_input = bc_pe_30_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_31_io_ve_input = bc_pe_15_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_31_io_input_valid = io_input_valid_31; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_31_io_iormac = io_iormac_31; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_32_clock = clock;
  assign bc_pe_32_reset = reset;
  assign bc_pe_32_io_ho_input = io_x_input_2; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_32_io_ve_input = bc_pe_16_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_32_io_input_valid = io_input_valid_32; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_32_io_iormac = io_iormac_32; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_33_clock = clock;
  assign bc_pe_33_reset = reset;
  assign bc_pe_33_io_ho_input = bc_pe_32_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_33_io_ve_input = bc_pe_17_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_33_io_input_valid = io_input_valid_33; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_33_io_iormac = io_iormac_33; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_34_clock = clock;
  assign bc_pe_34_reset = reset;
  assign bc_pe_34_io_ho_input = bc_pe_33_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_34_io_ve_input = bc_pe_18_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_34_io_input_valid = io_input_valid_34; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_34_io_iormac = io_iormac_34; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_35_clock = clock;
  assign bc_pe_35_reset = reset;
  assign bc_pe_35_io_ho_input = bc_pe_34_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_35_io_ve_input = bc_pe_19_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_35_io_input_valid = io_input_valid_35; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_35_io_iormac = io_iormac_35; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_36_clock = clock;
  assign bc_pe_36_reset = reset;
  assign bc_pe_36_io_ho_input = bc_pe_35_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_36_io_ve_input = bc_pe_20_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_36_io_input_valid = io_input_valid_36; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_36_io_iormac = io_iormac_36; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_37_clock = clock;
  assign bc_pe_37_reset = reset;
  assign bc_pe_37_io_ho_input = bc_pe_36_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_37_io_ve_input = bc_pe_21_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_37_io_input_valid = io_input_valid_37; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_37_io_iormac = io_iormac_37; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_38_clock = clock;
  assign bc_pe_38_reset = reset;
  assign bc_pe_38_io_ho_input = bc_pe_37_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_38_io_ve_input = bc_pe_22_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_38_io_input_valid = io_input_valid_38; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_38_io_iormac = io_iormac_38; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_39_clock = clock;
  assign bc_pe_39_reset = reset;
  assign bc_pe_39_io_ho_input = bc_pe_38_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_39_io_ve_input = bc_pe_23_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_39_io_input_valid = io_input_valid_39; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_39_io_iormac = io_iormac_39; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_40_clock = clock;
  assign bc_pe_40_reset = reset;
  assign bc_pe_40_io_ho_input = bc_pe_39_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_40_io_ve_input = bc_pe_24_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_40_io_input_valid = io_input_valid_40; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_40_io_iormac = io_iormac_40; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_41_clock = clock;
  assign bc_pe_41_reset = reset;
  assign bc_pe_41_io_ho_input = bc_pe_40_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_41_io_ve_input = bc_pe_25_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_41_io_input_valid = io_input_valid_41; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_41_io_iormac = io_iormac_41; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_42_clock = clock;
  assign bc_pe_42_reset = reset;
  assign bc_pe_42_io_ho_input = bc_pe_41_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_42_io_ve_input = bc_pe_26_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_42_io_input_valid = io_input_valid_42; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_42_io_iormac = io_iormac_42; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_43_clock = clock;
  assign bc_pe_43_reset = reset;
  assign bc_pe_43_io_ho_input = bc_pe_42_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_43_io_ve_input = bc_pe_27_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_43_io_input_valid = io_input_valid_43; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_43_io_iormac = io_iormac_43; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_44_clock = clock;
  assign bc_pe_44_reset = reset;
  assign bc_pe_44_io_ho_input = bc_pe_43_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_44_io_ve_input = bc_pe_28_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_44_io_input_valid = io_input_valid_44; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_44_io_iormac = io_iormac_44; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_45_clock = clock;
  assign bc_pe_45_reset = reset;
  assign bc_pe_45_io_ho_input = bc_pe_44_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_45_io_ve_input = bc_pe_29_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_45_io_input_valid = io_input_valid_45; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_45_io_iormac = io_iormac_45; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_46_clock = clock;
  assign bc_pe_46_reset = reset;
  assign bc_pe_46_io_ho_input = bc_pe_45_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_46_io_ve_input = bc_pe_30_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_46_io_input_valid = io_input_valid_46; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_46_io_iormac = io_iormac_46; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_47_clock = clock;
  assign bc_pe_47_reset = reset;
  assign bc_pe_47_io_ho_input = bc_pe_46_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_47_io_ve_input = bc_pe_31_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_47_io_input_valid = io_input_valid_47; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_47_io_iormac = io_iormac_47; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_48_clock = clock;
  assign bc_pe_48_reset = reset;
  assign bc_pe_48_io_ho_input = io_x_input_3; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_48_io_ve_input = bc_pe_32_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_48_io_input_valid = io_input_valid_48; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_48_io_iormac = io_iormac_48; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_49_clock = clock;
  assign bc_pe_49_reset = reset;
  assign bc_pe_49_io_ho_input = bc_pe_48_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_49_io_ve_input = bc_pe_33_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_49_io_input_valid = io_input_valid_49; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_49_io_iormac = io_iormac_49; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_50_clock = clock;
  assign bc_pe_50_reset = reset;
  assign bc_pe_50_io_ho_input = bc_pe_49_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_50_io_ve_input = bc_pe_34_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_50_io_input_valid = io_input_valid_50; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_50_io_iormac = io_iormac_50; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_51_clock = clock;
  assign bc_pe_51_reset = reset;
  assign bc_pe_51_io_ho_input = bc_pe_50_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_51_io_ve_input = bc_pe_35_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_51_io_input_valid = io_input_valid_51; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_51_io_iormac = io_iormac_51; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_52_clock = clock;
  assign bc_pe_52_reset = reset;
  assign bc_pe_52_io_ho_input = bc_pe_51_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_52_io_ve_input = bc_pe_36_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_52_io_input_valid = io_input_valid_52; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_52_io_iormac = io_iormac_52; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_53_clock = clock;
  assign bc_pe_53_reset = reset;
  assign bc_pe_53_io_ho_input = bc_pe_52_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_53_io_ve_input = bc_pe_37_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_53_io_input_valid = io_input_valid_53; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_53_io_iormac = io_iormac_53; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_54_clock = clock;
  assign bc_pe_54_reset = reset;
  assign bc_pe_54_io_ho_input = bc_pe_53_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_54_io_ve_input = bc_pe_38_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_54_io_input_valid = io_input_valid_54; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_54_io_iormac = io_iormac_54; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_55_clock = clock;
  assign bc_pe_55_reset = reset;
  assign bc_pe_55_io_ho_input = bc_pe_54_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_55_io_ve_input = bc_pe_39_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_55_io_input_valid = io_input_valid_55; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_55_io_iormac = io_iormac_55; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_56_clock = clock;
  assign bc_pe_56_reset = reset;
  assign bc_pe_56_io_ho_input = bc_pe_55_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_56_io_ve_input = bc_pe_40_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_56_io_input_valid = io_input_valid_56; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_56_io_iormac = io_iormac_56; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_57_clock = clock;
  assign bc_pe_57_reset = reset;
  assign bc_pe_57_io_ho_input = bc_pe_56_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_57_io_ve_input = bc_pe_41_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_57_io_input_valid = io_input_valid_57; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_57_io_iormac = io_iormac_57; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_58_clock = clock;
  assign bc_pe_58_reset = reset;
  assign bc_pe_58_io_ho_input = bc_pe_57_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_58_io_ve_input = bc_pe_42_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_58_io_input_valid = io_input_valid_58; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_58_io_iormac = io_iormac_58; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_59_clock = clock;
  assign bc_pe_59_reset = reset;
  assign bc_pe_59_io_ho_input = bc_pe_58_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_59_io_ve_input = bc_pe_43_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_59_io_input_valid = io_input_valid_59; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_59_io_iormac = io_iormac_59; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_60_clock = clock;
  assign bc_pe_60_reset = reset;
  assign bc_pe_60_io_ho_input = bc_pe_59_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_60_io_ve_input = bc_pe_44_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_60_io_input_valid = io_input_valid_60; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_60_io_iormac = io_iormac_60; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_61_clock = clock;
  assign bc_pe_61_reset = reset;
  assign bc_pe_61_io_ho_input = bc_pe_60_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_61_io_ve_input = bc_pe_45_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_61_io_input_valid = io_input_valid_61; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_61_io_iormac = io_iormac_61; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_62_clock = clock;
  assign bc_pe_62_reset = reset;
  assign bc_pe_62_io_ho_input = bc_pe_61_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_62_io_ve_input = bc_pe_46_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_62_io_input_valid = io_input_valid_62; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_62_io_iormac = io_iormac_62; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_63_clock = clock;
  assign bc_pe_63_reset = reset;
  assign bc_pe_63_io_ho_input = bc_pe_62_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_63_io_ve_input = bc_pe_47_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_63_io_input_valid = io_input_valid_63; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_63_io_iormac = io_iormac_63; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_64_clock = clock;
  assign bc_pe_64_reset = reset;
  assign bc_pe_64_io_ho_input = io_x_input_4; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_64_io_ve_input = bc_pe_48_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_64_io_input_valid = io_input_valid_64; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_64_io_iormac = io_iormac_64; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_65_clock = clock;
  assign bc_pe_65_reset = reset;
  assign bc_pe_65_io_ho_input = bc_pe_64_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_65_io_ve_input = bc_pe_49_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_65_io_input_valid = io_input_valid_65; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_65_io_iormac = io_iormac_65; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_66_clock = clock;
  assign bc_pe_66_reset = reset;
  assign bc_pe_66_io_ho_input = bc_pe_65_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_66_io_ve_input = bc_pe_50_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_66_io_input_valid = io_input_valid_66; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_66_io_iormac = io_iormac_66; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_67_clock = clock;
  assign bc_pe_67_reset = reset;
  assign bc_pe_67_io_ho_input = bc_pe_66_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_67_io_ve_input = bc_pe_51_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_67_io_input_valid = io_input_valid_67; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_67_io_iormac = io_iormac_67; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_68_clock = clock;
  assign bc_pe_68_reset = reset;
  assign bc_pe_68_io_ho_input = bc_pe_67_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_68_io_ve_input = bc_pe_52_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_68_io_input_valid = io_input_valid_68; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_68_io_iormac = io_iormac_68; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_69_clock = clock;
  assign bc_pe_69_reset = reset;
  assign bc_pe_69_io_ho_input = bc_pe_68_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_69_io_ve_input = bc_pe_53_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_69_io_input_valid = io_input_valid_69; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_69_io_iormac = io_iormac_69; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_70_clock = clock;
  assign bc_pe_70_reset = reset;
  assign bc_pe_70_io_ho_input = bc_pe_69_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_70_io_ve_input = bc_pe_54_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_70_io_input_valid = io_input_valid_70; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_70_io_iormac = io_iormac_70; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_71_clock = clock;
  assign bc_pe_71_reset = reset;
  assign bc_pe_71_io_ho_input = bc_pe_70_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_71_io_ve_input = bc_pe_55_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_71_io_input_valid = io_input_valid_71; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_71_io_iormac = io_iormac_71; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_72_clock = clock;
  assign bc_pe_72_reset = reset;
  assign bc_pe_72_io_ho_input = bc_pe_71_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_72_io_ve_input = bc_pe_56_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_72_io_input_valid = io_input_valid_72; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_72_io_iormac = io_iormac_72; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_73_clock = clock;
  assign bc_pe_73_reset = reset;
  assign bc_pe_73_io_ho_input = bc_pe_72_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_73_io_ve_input = bc_pe_57_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_73_io_input_valid = io_input_valid_73; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_73_io_iormac = io_iormac_73; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_74_clock = clock;
  assign bc_pe_74_reset = reset;
  assign bc_pe_74_io_ho_input = bc_pe_73_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_74_io_ve_input = bc_pe_58_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_74_io_input_valid = io_input_valid_74; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_74_io_iormac = io_iormac_74; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_75_clock = clock;
  assign bc_pe_75_reset = reset;
  assign bc_pe_75_io_ho_input = bc_pe_74_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_75_io_ve_input = bc_pe_59_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_75_io_input_valid = io_input_valid_75; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_75_io_iormac = io_iormac_75; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_76_clock = clock;
  assign bc_pe_76_reset = reset;
  assign bc_pe_76_io_ho_input = bc_pe_75_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_76_io_ve_input = bc_pe_60_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_76_io_input_valid = io_input_valid_76; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_76_io_iormac = io_iormac_76; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_77_clock = clock;
  assign bc_pe_77_reset = reset;
  assign bc_pe_77_io_ho_input = bc_pe_76_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_77_io_ve_input = bc_pe_61_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_77_io_input_valid = io_input_valid_77; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_77_io_iormac = io_iormac_77; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_78_clock = clock;
  assign bc_pe_78_reset = reset;
  assign bc_pe_78_io_ho_input = bc_pe_77_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_78_io_ve_input = bc_pe_62_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_78_io_input_valid = io_input_valid_78; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_78_io_iormac = io_iormac_78; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_79_clock = clock;
  assign bc_pe_79_reset = reset;
  assign bc_pe_79_io_ho_input = bc_pe_78_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_79_io_ve_input = bc_pe_63_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_79_io_input_valid = io_input_valid_79; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_79_io_iormac = io_iormac_79; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_80_clock = clock;
  assign bc_pe_80_reset = reset;
  assign bc_pe_80_io_ho_input = io_x_input_5; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_80_io_ve_input = bc_pe_64_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_80_io_input_valid = io_input_valid_80; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_80_io_iormac = io_iormac_80; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_81_clock = clock;
  assign bc_pe_81_reset = reset;
  assign bc_pe_81_io_ho_input = bc_pe_80_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_81_io_ve_input = bc_pe_65_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_81_io_input_valid = io_input_valid_81; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_81_io_iormac = io_iormac_81; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_82_clock = clock;
  assign bc_pe_82_reset = reset;
  assign bc_pe_82_io_ho_input = bc_pe_81_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_82_io_ve_input = bc_pe_66_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_82_io_input_valid = io_input_valid_82; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_82_io_iormac = io_iormac_82; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_83_clock = clock;
  assign bc_pe_83_reset = reset;
  assign bc_pe_83_io_ho_input = bc_pe_82_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_83_io_ve_input = bc_pe_67_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_83_io_input_valid = io_input_valid_83; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_83_io_iormac = io_iormac_83; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_84_clock = clock;
  assign bc_pe_84_reset = reset;
  assign bc_pe_84_io_ho_input = bc_pe_83_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_84_io_ve_input = bc_pe_68_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_84_io_input_valid = io_input_valid_84; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_84_io_iormac = io_iormac_84; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_85_clock = clock;
  assign bc_pe_85_reset = reset;
  assign bc_pe_85_io_ho_input = bc_pe_84_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_85_io_ve_input = bc_pe_69_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_85_io_input_valid = io_input_valid_85; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_85_io_iormac = io_iormac_85; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_86_clock = clock;
  assign bc_pe_86_reset = reset;
  assign bc_pe_86_io_ho_input = bc_pe_85_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_86_io_ve_input = bc_pe_70_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_86_io_input_valid = io_input_valid_86; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_86_io_iormac = io_iormac_86; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_87_clock = clock;
  assign bc_pe_87_reset = reset;
  assign bc_pe_87_io_ho_input = bc_pe_86_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_87_io_ve_input = bc_pe_71_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_87_io_input_valid = io_input_valid_87; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_87_io_iormac = io_iormac_87; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_88_clock = clock;
  assign bc_pe_88_reset = reset;
  assign bc_pe_88_io_ho_input = bc_pe_87_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_88_io_ve_input = bc_pe_72_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_88_io_input_valid = io_input_valid_88; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_88_io_iormac = io_iormac_88; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_89_clock = clock;
  assign bc_pe_89_reset = reset;
  assign bc_pe_89_io_ho_input = bc_pe_88_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_89_io_ve_input = bc_pe_73_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_89_io_input_valid = io_input_valid_89; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_89_io_iormac = io_iormac_89; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_90_clock = clock;
  assign bc_pe_90_reset = reset;
  assign bc_pe_90_io_ho_input = bc_pe_89_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_90_io_ve_input = bc_pe_74_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_90_io_input_valid = io_input_valid_90; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_90_io_iormac = io_iormac_90; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_91_clock = clock;
  assign bc_pe_91_reset = reset;
  assign bc_pe_91_io_ho_input = bc_pe_90_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_91_io_ve_input = bc_pe_75_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_91_io_input_valid = io_input_valid_91; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_91_io_iormac = io_iormac_91; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_92_clock = clock;
  assign bc_pe_92_reset = reset;
  assign bc_pe_92_io_ho_input = bc_pe_91_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_92_io_ve_input = bc_pe_76_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_92_io_input_valid = io_input_valid_92; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_92_io_iormac = io_iormac_92; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_93_clock = clock;
  assign bc_pe_93_reset = reset;
  assign bc_pe_93_io_ho_input = bc_pe_92_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_93_io_ve_input = bc_pe_77_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_93_io_input_valid = io_input_valid_93; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_93_io_iormac = io_iormac_93; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_94_clock = clock;
  assign bc_pe_94_reset = reset;
  assign bc_pe_94_io_ho_input = bc_pe_93_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_94_io_ve_input = bc_pe_78_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_94_io_input_valid = io_input_valid_94; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_94_io_iormac = io_iormac_94; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_95_clock = clock;
  assign bc_pe_95_reset = reset;
  assign bc_pe_95_io_ho_input = bc_pe_94_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_95_io_ve_input = bc_pe_79_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_95_io_input_valid = io_input_valid_95; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_95_io_iormac = io_iormac_95; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_96_clock = clock;
  assign bc_pe_96_reset = reset;
  assign bc_pe_96_io_ho_input = io_x_input_6; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_96_io_ve_input = bc_pe_80_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_96_io_input_valid = io_input_valid_96; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_96_io_iormac = io_iormac_96; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_97_clock = clock;
  assign bc_pe_97_reset = reset;
  assign bc_pe_97_io_ho_input = bc_pe_96_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_97_io_ve_input = bc_pe_81_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_97_io_input_valid = io_input_valid_97; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_97_io_iormac = io_iormac_97; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_98_clock = clock;
  assign bc_pe_98_reset = reset;
  assign bc_pe_98_io_ho_input = bc_pe_97_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_98_io_ve_input = bc_pe_82_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_98_io_input_valid = io_input_valid_98; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_98_io_iormac = io_iormac_98; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_99_clock = clock;
  assign bc_pe_99_reset = reset;
  assign bc_pe_99_io_ho_input = bc_pe_98_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_99_io_ve_input = bc_pe_83_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_99_io_input_valid = io_input_valid_99; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_99_io_iormac = io_iormac_99; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_100_clock = clock;
  assign bc_pe_100_reset = reset;
  assign bc_pe_100_io_ho_input = bc_pe_99_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_100_io_ve_input = bc_pe_84_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_100_io_input_valid = io_input_valid_100; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_100_io_iormac = io_iormac_100; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_101_clock = clock;
  assign bc_pe_101_reset = reset;
  assign bc_pe_101_io_ho_input = bc_pe_100_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_101_io_ve_input = bc_pe_85_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_101_io_input_valid = io_input_valid_101; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_101_io_iormac = io_iormac_101; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_102_clock = clock;
  assign bc_pe_102_reset = reset;
  assign bc_pe_102_io_ho_input = bc_pe_101_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_102_io_ve_input = bc_pe_86_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_102_io_input_valid = io_input_valid_102; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_102_io_iormac = io_iormac_102; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_103_clock = clock;
  assign bc_pe_103_reset = reset;
  assign bc_pe_103_io_ho_input = bc_pe_102_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_103_io_ve_input = bc_pe_87_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_103_io_input_valid = io_input_valid_103; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_103_io_iormac = io_iormac_103; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_104_clock = clock;
  assign bc_pe_104_reset = reset;
  assign bc_pe_104_io_ho_input = bc_pe_103_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_104_io_ve_input = bc_pe_88_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_104_io_input_valid = io_input_valid_104; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_104_io_iormac = io_iormac_104; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_105_clock = clock;
  assign bc_pe_105_reset = reset;
  assign bc_pe_105_io_ho_input = bc_pe_104_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_105_io_ve_input = bc_pe_89_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_105_io_input_valid = io_input_valid_105; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_105_io_iormac = io_iormac_105; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_106_clock = clock;
  assign bc_pe_106_reset = reset;
  assign bc_pe_106_io_ho_input = bc_pe_105_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_106_io_ve_input = bc_pe_90_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_106_io_input_valid = io_input_valid_106; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_106_io_iormac = io_iormac_106; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_107_clock = clock;
  assign bc_pe_107_reset = reset;
  assign bc_pe_107_io_ho_input = bc_pe_106_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_107_io_ve_input = bc_pe_91_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_107_io_input_valid = io_input_valid_107; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_107_io_iormac = io_iormac_107; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_108_clock = clock;
  assign bc_pe_108_reset = reset;
  assign bc_pe_108_io_ho_input = bc_pe_107_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_108_io_ve_input = bc_pe_92_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_108_io_input_valid = io_input_valid_108; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_108_io_iormac = io_iormac_108; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_109_clock = clock;
  assign bc_pe_109_reset = reset;
  assign bc_pe_109_io_ho_input = bc_pe_108_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_109_io_ve_input = bc_pe_93_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_109_io_input_valid = io_input_valid_109; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_109_io_iormac = io_iormac_109; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_110_clock = clock;
  assign bc_pe_110_reset = reset;
  assign bc_pe_110_io_ho_input = bc_pe_109_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_110_io_ve_input = bc_pe_94_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_110_io_input_valid = io_input_valid_110; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_110_io_iormac = io_iormac_110; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_111_clock = clock;
  assign bc_pe_111_reset = reset;
  assign bc_pe_111_io_ho_input = bc_pe_110_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_111_io_ve_input = bc_pe_95_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_111_io_input_valid = io_input_valid_111; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_111_io_iormac = io_iormac_111; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_112_clock = clock;
  assign bc_pe_112_reset = reset;
  assign bc_pe_112_io_ho_input = io_x_input_7; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_112_io_ve_input = bc_pe_96_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_112_io_input_valid = io_input_valid_112; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_112_io_iormac = io_iormac_112; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_113_clock = clock;
  assign bc_pe_113_reset = reset;
  assign bc_pe_113_io_ho_input = bc_pe_112_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_113_io_ve_input = bc_pe_97_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_113_io_input_valid = io_input_valid_113; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_113_io_iormac = io_iormac_113; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_114_clock = clock;
  assign bc_pe_114_reset = reset;
  assign bc_pe_114_io_ho_input = bc_pe_113_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_114_io_ve_input = bc_pe_98_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_114_io_input_valid = io_input_valid_114; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_114_io_iormac = io_iormac_114; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_115_clock = clock;
  assign bc_pe_115_reset = reset;
  assign bc_pe_115_io_ho_input = bc_pe_114_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_115_io_ve_input = bc_pe_99_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_115_io_input_valid = io_input_valid_115; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_115_io_iormac = io_iormac_115; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_116_clock = clock;
  assign bc_pe_116_reset = reset;
  assign bc_pe_116_io_ho_input = bc_pe_115_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_116_io_ve_input = bc_pe_100_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_116_io_input_valid = io_input_valid_116; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_116_io_iormac = io_iormac_116; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_117_clock = clock;
  assign bc_pe_117_reset = reset;
  assign bc_pe_117_io_ho_input = bc_pe_116_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_117_io_ve_input = bc_pe_101_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_117_io_input_valid = io_input_valid_117; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_117_io_iormac = io_iormac_117; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_118_clock = clock;
  assign bc_pe_118_reset = reset;
  assign bc_pe_118_io_ho_input = bc_pe_117_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_118_io_ve_input = bc_pe_102_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_118_io_input_valid = io_input_valid_118; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_118_io_iormac = io_iormac_118; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_119_clock = clock;
  assign bc_pe_119_reset = reset;
  assign bc_pe_119_io_ho_input = bc_pe_118_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_119_io_ve_input = bc_pe_103_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_119_io_input_valid = io_input_valid_119; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_119_io_iormac = io_iormac_119; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_120_clock = clock;
  assign bc_pe_120_reset = reset;
  assign bc_pe_120_io_ho_input = bc_pe_119_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_120_io_ve_input = bc_pe_104_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_120_io_input_valid = io_input_valid_120; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_120_io_iormac = io_iormac_120; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_121_clock = clock;
  assign bc_pe_121_reset = reset;
  assign bc_pe_121_io_ho_input = bc_pe_120_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_121_io_ve_input = bc_pe_105_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_121_io_input_valid = io_input_valid_121; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_121_io_iormac = io_iormac_121; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_122_clock = clock;
  assign bc_pe_122_reset = reset;
  assign bc_pe_122_io_ho_input = bc_pe_121_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_122_io_ve_input = bc_pe_106_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_122_io_input_valid = io_input_valid_122; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_122_io_iormac = io_iormac_122; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_123_clock = clock;
  assign bc_pe_123_reset = reset;
  assign bc_pe_123_io_ho_input = bc_pe_122_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_123_io_ve_input = bc_pe_107_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_123_io_input_valid = io_input_valid_123; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_123_io_iormac = io_iormac_123; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_124_clock = clock;
  assign bc_pe_124_reset = reset;
  assign bc_pe_124_io_ho_input = bc_pe_123_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_124_io_ve_input = bc_pe_108_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_124_io_input_valid = io_input_valid_124; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_124_io_iormac = io_iormac_124; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_125_clock = clock;
  assign bc_pe_125_reset = reset;
  assign bc_pe_125_io_ho_input = bc_pe_124_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_125_io_ve_input = bc_pe_109_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_125_io_input_valid = io_input_valid_125; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_125_io_iormac = io_iormac_125; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_126_clock = clock;
  assign bc_pe_126_reset = reset;
  assign bc_pe_126_io_ho_input = bc_pe_125_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_126_io_ve_input = bc_pe_110_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_126_io_input_valid = io_input_valid_126; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_126_io_iormac = io_iormac_126; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_127_clock = clock;
  assign bc_pe_127_reset = reset;
  assign bc_pe_127_io_ho_input = bc_pe_126_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_127_io_ve_input = bc_pe_111_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_127_io_input_valid = io_input_valid_127; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_127_io_iormac = io_iormac_127; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_128_clock = clock;
  assign bc_pe_128_reset = reset;
  assign bc_pe_128_io_ho_input = io_x_input_8; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_128_io_ve_input = bc_pe_112_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_128_io_input_valid = io_input_valid_128; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_128_io_iormac = io_iormac_128; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_129_clock = clock;
  assign bc_pe_129_reset = reset;
  assign bc_pe_129_io_ho_input = bc_pe_128_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_129_io_ve_input = bc_pe_113_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_129_io_input_valid = io_input_valid_129; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_129_io_iormac = io_iormac_129; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_130_clock = clock;
  assign bc_pe_130_reset = reset;
  assign bc_pe_130_io_ho_input = bc_pe_129_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_130_io_ve_input = bc_pe_114_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_130_io_input_valid = io_input_valid_130; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_130_io_iormac = io_iormac_130; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_131_clock = clock;
  assign bc_pe_131_reset = reset;
  assign bc_pe_131_io_ho_input = bc_pe_130_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_131_io_ve_input = bc_pe_115_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_131_io_input_valid = io_input_valid_131; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_131_io_iormac = io_iormac_131; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_132_clock = clock;
  assign bc_pe_132_reset = reset;
  assign bc_pe_132_io_ho_input = bc_pe_131_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_132_io_ve_input = bc_pe_116_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_132_io_input_valid = io_input_valid_132; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_132_io_iormac = io_iormac_132; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_133_clock = clock;
  assign bc_pe_133_reset = reset;
  assign bc_pe_133_io_ho_input = bc_pe_132_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_133_io_ve_input = bc_pe_117_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_133_io_input_valid = io_input_valid_133; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_133_io_iormac = io_iormac_133; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_134_clock = clock;
  assign bc_pe_134_reset = reset;
  assign bc_pe_134_io_ho_input = bc_pe_133_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_134_io_ve_input = bc_pe_118_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_134_io_input_valid = io_input_valid_134; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_134_io_iormac = io_iormac_134; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_135_clock = clock;
  assign bc_pe_135_reset = reset;
  assign bc_pe_135_io_ho_input = bc_pe_134_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_135_io_ve_input = bc_pe_119_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_135_io_input_valid = io_input_valid_135; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_135_io_iormac = io_iormac_135; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_136_clock = clock;
  assign bc_pe_136_reset = reset;
  assign bc_pe_136_io_ho_input = bc_pe_135_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_136_io_ve_input = bc_pe_120_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_136_io_input_valid = io_input_valid_136; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_136_io_iormac = io_iormac_136; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_137_clock = clock;
  assign bc_pe_137_reset = reset;
  assign bc_pe_137_io_ho_input = bc_pe_136_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_137_io_ve_input = bc_pe_121_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_137_io_input_valid = io_input_valid_137; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_137_io_iormac = io_iormac_137; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_138_clock = clock;
  assign bc_pe_138_reset = reset;
  assign bc_pe_138_io_ho_input = bc_pe_137_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_138_io_ve_input = bc_pe_122_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_138_io_input_valid = io_input_valid_138; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_138_io_iormac = io_iormac_138; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_139_clock = clock;
  assign bc_pe_139_reset = reset;
  assign bc_pe_139_io_ho_input = bc_pe_138_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_139_io_ve_input = bc_pe_123_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_139_io_input_valid = io_input_valid_139; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_139_io_iormac = io_iormac_139; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_140_clock = clock;
  assign bc_pe_140_reset = reset;
  assign bc_pe_140_io_ho_input = bc_pe_139_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_140_io_ve_input = bc_pe_124_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_140_io_input_valid = io_input_valid_140; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_140_io_iormac = io_iormac_140; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_141_clock = clock;
  assign bc_pe_141_reset = reset;
  assign bc_pe_141_io_ho_input = bc_pe_140_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_141_io_ve_input = bc_pe_125_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_141_io_input_valid = io_input_valid_141; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_141_io_iormac = io_iormac_141; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_142_clock = clock;
  assign bc_pe_142_reset = reset;
  assign bc_pe_142_io_ho_input = bc_pe_141_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_142_io_ve_input = bc_pe_126_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_142_io_input_valid = io_input_valid_142; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_142_io_iormac = io_iormac_142; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_143_clock = clock;
  assign bc_pe_143_reset = reset;
  assign bc_pe_143_io_ho_input = bc_pe_142_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_143_io_ve_input = bc_pe_127_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_143_io_input_valid = io_input_valid_143; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_143_io_iormac = io_iormac_143; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_144_clock = clock;
  assign bc_pe_144_reset = reset;
  assign bc_pe_144_io_ho_input = io_x_input_9; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_144_io_ve_input = bc_pe_128_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_144_io_input_valid = io_input_valid_144; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_144_io_iormac = io_iormac_144; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_145_clock = clock;
  assign bc_pe_145_reset = reset;
  assign bc_pe_145_io_ho_input = bc_pe_144_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_145_io_ve_input = bc_pe_129_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_145_io_input_valid = io_input_valid_145; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_145_io_iormac = io_iormac_145; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_146_clock = clock;
  assign bc_pe_146_reset = reset;
  assign bc_pe_146_io_ho_input = bc_pe_145_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_146_io_ve_input = bc_pe_130_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_146_io_input_valid = io_input_valid_146; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_146_io_iormac = io_iormac_146; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_147_clock = clock;
  assign bc_pe_147_reset = reset;
  assign bc_pe_147_io_ho_input = bc_pe_146_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_147_io_ve_input = bc_pe_131_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_147_io_input_valid = io_input_valid_147; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_147_io_iormac = io_iormac_147; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_148_clock = clock;
  assign bc_pe_148_reset = reset;
  assign bc_pe_148_io_ho_input = bc_pe_147_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_148_io_ve_input = bc_pe_132_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_148_io_input_valid = io_input_valid_148; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_148_io_iormac = io_iormac_148; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_149_clock = clock;
  assign bc_pe_149_reset = reset;
  assign bc_pe_149_io_ho_input = bc_pe_148_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_149_io_ve_input = bc_pe_133_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_149_io_input_valid = io_input_valid_149; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_149_io_iormac = io_iormac_149; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_150_clock = clock;
  assign bc_pe_150_reset = reset;
  assign bc_pe_150_io_ho_input = bc_pe_149_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_150_io_ve_input = bc_pe_134_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_150_io_input_valid = io_input_valid_150; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_150_io_iormac = io_iormac_150; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_151_clock = clock;
  assign bc_pe_151_reset = reset;
  assign bc_pe_151_io_ho_input = bc_pe_150_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_151_io_ve_input = bc_pe_135_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_151_io_input_valid = io_input_valid_151; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_151_io_iormac = io_iormac_151; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_152_clock = clock;
  assign bc_pe_152_reset = reset;
  assign bc_pe_152_io_ho_input = bc_pe_151_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_152_io_ve_input = bc_pe_136_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_152_io_input_valid = io_input_valid_152; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_152_io_iormac = io_iormac_152; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_153_clock = clock;
  assign bc_pe_153_reset = reset;
  assign bc_pe_153_io_ho_input = bc_pe_152_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_153_io_ve_input = bc_pe_137_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_153_io_input_valid = io_input_valid_153; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_153_io_iormac = io_iormac_153; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_154_clock = clock;
  assign bc_pe_154_reset = reset;
  assign bc_pe_154_io_ho_input = bc_pe_153_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_154_io_ve_input = bc_pe_138_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_154_io_input_valid = io_input_valid_154; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_154_io_iormac = io_iormac_154; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_155_clock = clock;
  assign bc_pe_155_reset = reset;
  assign bc_pe_155_io_ho_input = bc_pe_154_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_155_io_ve_input = bc_pe_139_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_155_io_input_valid = io_input_valid_155; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_155_io_iormac = io_iormac_155; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_156_clock = clock;
  assign bc_pe_156_reset = reset;
  assign bc_pe_156_io_ho_input = bc_pe_155_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_156_io_ve_input = bc_pe_140_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_156_io_input_valid = io_input_valid_156; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_156_io_iormac = io_iormac_156; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_157_clock = clock;
  assign bc_pe_157_reset = reset;
  assign bc_pe_157_io_ho_input = bc_pe_156_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_157_io_ve_input = bc_pe_141_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_157_io_input_valid = io_input_valid_157; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_157_io_iormac = io_iormac_157; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_158_clock = clock;
  assign bc_pe_158_reset = reset;
  assign bc_pe_158_io_ho_input = bc_pe_157_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_158_io_ve_input = bc_pe_142_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_158_io_input_valid = io_input_valid_158; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_158_io_iormac = io_iormac_158; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_159_clock = clock;
  assign bc_pe_159_reset = reset;
  assign bc_pe_159_io_ho_input = bc_pe_158_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_159_io_ve_input = bc_pe_143_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_159_io_input_valid = io_input_valid_159; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_159_io_iormac = io_iormac_159; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_160_clock = clock;
  assign bc_pe_160_reset = reset;
  assign bc_pe_160_io_ho_input = io_x_input_10; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_160_io_ve_input = bc_pe_144_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_160_io_input_valid = io_input_valid_160; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_160_io_iormac = io_iormac_160; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_161_clock = clock;
  assign bc_pe_161_reset = reset;
  assign bc_pe_161_io_ho_input = bc_pe_160_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_161_io_ve_input = bc_pe_145_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_161_io_input_valid = io_input_valid_161; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_161_io_iormac = io_iormac_161; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_162_clock = clock;
  assign bc_pe_162_reset = reset;
  assign bc_pe_162_io_ho_input = bc_pe_161_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_162_io_ve_input = bc_pe_146_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_162_io_input_valid = io_input_valid_162; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_162_io_iormac = io_iormac_162; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_163_clock = clock;
  assign bc_pe_163_reset = reset;
  assign bc_pe_163_io_ho_input = bc_pe_162_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_163_io_ve_input = bc_pe_147_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_163_io_input_valid = io_input_valid_163; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_163_io_iormac = io_iormac_163; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_164_clock = clock;
  assign bc_pe_164_reset = reset;
  assign bc_pe_164_io_ho_input = bc_pe_163_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_164_io_ve_input = bc_pe_148_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_164_io_input_valid = io_input_valid_164; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_164_io_iormac = io_iormac_164; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_165_clock = clock;
  assign bc_pe_165_reset = reset;
  assign bc_pe_165_io_ho_input = bc_pe_164_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_165_io_ve_input = bc_pe_149_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_165_io_input_valid = io_input_valid_165; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_165_io_iormac = io_iormac_165; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_166_clock = clock;
  assign bc_pe_166_reset = reset;
  assign bc_pe_166_io_ho_input = bc_pe_165_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_166_io_ve_input = bc_pe_150_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_166_io_input_valid = io_input_valid_166; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_166_io_iormac = io_iormac_166; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_167_clock = clock;
  assign bc_pe_167_reset = reset;
  assign bc_pe_167_io_ho_input = bc_pe_166_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_167_io_ve_input = bc_pe_151_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_167_io_input_valid = io_input_valid_167; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_167_io_iormac = io_iormac_167; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_168_clock = clock;
  assign bc_pe_168_reset = reset;
  assign bc_pe_168_io_ho_input = bc_pe_167_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_168_io_ve_input = bc_pe_152_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_168_io_input_valid = io_input_valid_168; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_168_io_iormac = io_iormac_168; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_169_clock = clock;
  assign bc_pe_169_reset = reset;
  assign bc_pe_169_io_ho_input = bc_pe_168_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_169_io_ve_input = bc_pe_153_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_169_io_input_valid = io_input_valid_169; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_169_io_iormac = io_iormac_169; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_170_clock = clock;
  assign bc_pe_170_reset = reset;
  assign bc_pe_170_io_ho_input = bc_pe_169_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_170_io_ve_input = bc_pe_154_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_170_io_input_valid = io_input_valid_170; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_170_io_iormac = io_iormac_170; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_171_clock = clock;
  assign bc_pe_171_reset = reset;
  assign bc_pe_171_io_ho_input = bc_pe_170_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_171_io_ve_input = bc_pe_155_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_171_io_input_valid = io_input_valid_171; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_171_io_iormac = io_iormac_171; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_172_clock = clock;
  assign bc_pe_172_reset = reset;
  assign bc_pe_172_io_ho_input = bc_pe_171_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_172_io_ve_input = bc_pe_156_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_172_io_input_valid = io_input_valid_172; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_172_io_iormac = io_iormac_172; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_173_clock = clock;
  assign bc_pe_173_reset = reset;
  assign bc_pe_173_io_ho_input = bc_pe_172_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_173_io_ve_input = bc_pe_157_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_173_io_input_valid = io_input_valid_173; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_173_io_iormac = io_iormac_173; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_174_clock = clock;
  assign bc_pe_174_reset = reset;
  assign bc_pe_174_io_ho_input = bc_pe_173_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_174_io_ve_input = bc_pe_158_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_174_io_input_valid = io_input_valid_174; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_174_io_iormac = io_iormac_174; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_175_clock = clock;
  assign bc_pe_175_reset = reset;
  assign bc_pe_175_io_ho_input = bc_pe_174_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_175_io_ve_input = bc_pe_159_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_175_io_input_valid = io_input_valid_175; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_175_io_iormac = io_iormac_175; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_176_clock = clock;
  assign bc_pe_176_reset = reset;
  assign bc_pe_176_io_ho_input = io_x_input_11; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_176_io_ve_input = bc_pe_160_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_176_io_input_valid = io_input_valid_176; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_176_io_iormac = io_iormac_176; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_177_clock = clock;
  assign bc_pe_177_reset = reset;
  assign bc_pe_177_io_ho_input = bc_pe_176_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_177_io_ve_input = bc_pe_161_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_177_io_input_valid = io_input_valid_177; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_177_io_iormac = io_iormac_177; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_178_clock = clock;
  assign bc_pe_178_reset = reset;
  assign bc_pe_178_io_ho_input = bc_pe_177_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_178_io_ve_input = bc_pe_162_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_178_io_input_valid = io_input_valid_178; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_178_io_iormac = io_iormac_178; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_179_clock = clock;
  assign bc_pe_179_reset = reset;
  assign bc_pe_179_io_ho_input = bc_pe_178_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_179_io_ve_input = bc_pe_163_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_179_io_input_valid = io_input_valid_179; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_179_io_iormac = io_iormac_179; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_180_clock = clock;
  assign bc_pe_180_reset = reset;
  assign bc_pe_180_io_ho_input = bc_pe_179_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_180_io_ve_input = bc_pe_164_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_180_io_input_valid = io_input_valid_180; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_180_io_iormac = io_iormac_180; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_181_clock = clock;
  assign bc_pe_181_reset = reset;
  assign bc_pe_181_io_ho_input = bc_pe_180_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_181_io_ve_input = bc_pe_165_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_181_io_input_valid = io_input_valid_181; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_181_io_iormac = io_iormac_181; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_182_clock = clock;
  assign bc_pe_182_reset = reset;
  assign bc_pe_182_io_ho_input = bc_pe_181_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_182_io_ve_input = bc_pe_166_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_182_io_input_valid = io_input_valid_182; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_182_io_iormac = io_iormac_182; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_183_clock = clock;
  assign bc_pe_183_reset = reset;
  assign bc_pe_183_io_ho_input = bc_pe_182_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_183_io_ve_input = bc_pe_167_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_183_io_input_valid = io_input_valid_183; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_183_io_iormac = io_iormac_183; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_184_clock = clock;
  assign bc_pe_184_reset = reset;
  assign bc_pe_184_io_ho_input = bc_pe_183_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_184_io_ve_input = bc_pe_168_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_184_io_input_valid = io_input_valid_184; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_184_io_iormac = io_iormac_184; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_185_clock = clock;
  assign bc_pe_185_reset = reset;
  assign bc_pe_185_io_ho_input = bc_pe_184_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_185_io_ve_input = bc_pe_169_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_185_io_input_valid = io_input_valid_185; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_185_io_iormac = io_iormac_185; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_186_clock = clock;
  assign bc_pe_186_reset = reset;
  assign bc_pe_186_io_ho_input = bc_pe_185_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_186_io_ve_input = bc_pe_170_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_186_io_input_valid = io_input_valid_186; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_186_io_iormac = io_iormac_186; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_187_clock = clock;
  assign bc_pe_187_reset = reset;
  assign bc_pe_187_io_ho_input = bc_pe_186_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_187_io_ve_input = bc_pe_171_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_187_io_input_valid = io_input_valid_187; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_187_io_iormac = io_iormac_187; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_188_clock = clock;
  assign bc_pe_188_reset = reset;
  assign bc_pe_188_io_ho_input = bc_pe_187_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_188_io_ve_input = bc_pe_172_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_188_io_input_valid = io_input_valid_188; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_188_io_iormac = io_iormac_188; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_189_clock = clock;
  assign bc_pe_189_reset = reset;
  assign bc_pe_189_io_ho_input = bc_pe_188_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_189_io_ve_input = bc_pe_173_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_189_io_input_valid = io_input_valid_189; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_189_io_iormac = io_iormac_189; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_190_clock = clock;
  assign bc_pe_190_reset = reset;
  assign bc_pe_190_io_ho_input = bc_pe_189_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_190_io_ve_input = bc_pe_174_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_190_io_input_valid = io_input_valid_190; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_190_io_iormac = io_iormac_190; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_191_clock = clock;
  assign bc_pe_191_reset = reset;
  assign bc_pe_191_io_ho_input = bc_pe_190_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_191_io_ve_input = bc_pe_175_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_191_io_input_valid = io_input_valid_191; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_191_io_iormac = io_iormac_191; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_192_clock = clock;
  assign bc_pe_192_reset = reset;
  assign bc_pe_192_io_ho_input = io_x_input_12; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_192_io_ve_input = bc_pe_176_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_192_io_input_valid = io_input_valid_192; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_192_io_iormac = io_iormac_192; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_193_clock = clock;
  assign bc_pe_193_reset = reset;
  assign bc_pe_193_io_ho_input = bc_pe_192_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_193_io_ve_input = bc_pe_177_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_193_io_input_valid = io_input_valid_193; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_193_io_iormac = io_iormac_193; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_194_clock = clock;
  assign bc_pe_194_reset = reset;
  assign bc_pe_194_io_ho_input = bc_pe_193_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_194_io_ve_input = bc_pe_178_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_194_io_input_valid = io_input_valid_194; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_194_io_iormac = io_iormac_194; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_195_clock = clock;
  assign bc_pe_195_reset = reset;
  assign bc_pe_195_io_ho_input = bc_pe_194_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_195_io_ve_input = bc_pe_179_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_195_io_input_valid = io_input_valid_195; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_195_io_iormac = io_iormac_195; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_196_clock = clock;
  assign bc_pe_196_reset = reset;
  assign bc_pe_196_io_ho_input = bc_pe_195_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_196_io_ve_input = bc_pe_180_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_196_io_input_valid = io_input_valid_196; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_196_io_iormac = io_iormac_196; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_197_clock = clock;
  assign bc_pe_197_reset = reset;
  assign bc_pe_197_io_ho_input = bc_pe_196_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_197_io_ve_input = bc_pe_181_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_197_io_input_valid = io_input_valid_197; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_197_io_iormac = io_iormac_197; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_198_clock = clock;
  assign bc_pe_198_reset = reset;
  assign bc_pe_198_io_ho_input = bc_pe_197_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_198_io_ve_input = bc_pe_182_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_198_io_input_valid = io_input_valid_198; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_198_io_iormac = io_iormac_198; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_199_clock = clock;
  assign bc_pe_199_reset = reset;
  assign bc_pe_199_io_ho_input = bc_pe_198_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_199_io_ve_input = bc_pe_183_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_199_io_input_valid = io_input_valid_199; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_199_io_iormac = io_iormac_199; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_200_clock = clock;
  assign bc_pe_200_reset = reset;
  assign bc_pe_200_io_ho_input = bc_pe_199_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_200_io_ve_input = bc_pe_184_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_200_io_input_valid = io_input_valid_200; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_200_io_iormac = io_iormac_200; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_201_clock = clock;
  assign bc_pe_201_reset = reset;
  assign bc_pe_201_io_ho_input = bc_pe_200_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_201_io_ve_input = bc_pe_185_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_201_io_input_valid = io_input_valid_201; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_201_io_iormac = io_iormac_201; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_202_clock = clock;
  assign bc_pe_202_reset = reset;
  assign bc_pe_202_io_ho_input = bc_pe_201_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_202_io_ve_input = bc_pe_186_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_202_io_input_valid = io_input_valid_202; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_202_io_iormac = io_iormac_202; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_203_clock = clock;
  assign bc_pe_203_reset = reset;
  assign bc_pe_203_io_ho_input = bc_pe_202_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_203_io_ve_input = bc_pe_187_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_203_io_input_valid = io_input_valid_203; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_203_io_iormac = io_iormac_203; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_204_clock = clock;
  assign bc_pe_204_reset = reset;
  assign bc_pe_204_io_ho_input = bc_pe_203_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_204_io_ve_input = bc_pe_188_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_204_io_input_valid = io_input_valid_204; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_204_io_iormac = io_iormac_204; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_205_clock = clock;
  assign bc_pe_205_reset = reset;
  assign bc_pe_205_io_ho_input = bc_pe_204_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_205_io_ve_input = bc_pe_189_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_205_io_input_valid = io_input_valid_205; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_205_io_iormac = io_iormac_205; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_206_clock = clock;
  assign bc_pe_206_reset = reset;
  assign bc_pe_206_io_ho_input = bc_pe_205_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_206_io_ve_input = bc_pe_190_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_206_io_input_valid = io_input_valid_206; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_206_io_iormac = io_iormac_206; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_207_clock = clock;
  assign bc_pe_207_reset = reset;
  assign bc_pe_207_io_ho_input = bc_pe_206_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_207_io_ve_input = bc_pe_191_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_207_io_input_valid = io_input_valid_207; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_207_io_iormac = io_iormac_207; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_208_clock = clock;
  assign bc_pe_208_reset = reset;
  assign bc_pe_208_io_ho_input = io_x_input_13; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_208_io_ve_input = bc_pe_192_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_208_io_input_valid = io_input_valid_208; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_208_io_iormac = io_iormac_208; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_209_clock = clock;
  assign bc_pe_209_reset = reset;
  assign bc_pe_209_io_ho_input = bc_pe_208_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_209_io_ve_input = bc_pe_193_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_209_io_input_valid = io_input_valid_209; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_209_io_iormac = io_iormac_209; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_210_clock = clock;
  assign bc_pe_210_reset = reset;
  assign bc_pe_210_io_ho_input = bc_pe_209_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_210_io_ve_input = bc_pe_194_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_210_io_input_valid = io_input_valid_210; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_210_io_iormac = io_iormac_210; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_211_clock = clock;
  assign bc_pe_211_reset = reset;
  assign bc_pe_211_io_ho_input = bc_pe_210_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_211_io_ve_input = bc_pe_195_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_211_io_input_valid = io_input_valid_211; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_211_io_iormac = io_iormac_211; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_212_clock = clock;
  assign bc_pe_212_reset = reset;
  assign bc_pe_212_io_ho_input = bc_pe_211_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_212_io_ve_input = bc_pe_196_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_212_io_input_valid = io_input_valid_212; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_212_io_iormac = io_iormac_212; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_213_clock = clock;
  assign bc_pe_213_reset = reset;
  assign bc_pe_213_io_ho_input = bc_pe_212_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_213_io_ve_input = bc_pe_197_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_213_io_input_valid = io_input_valid_213; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_213_io_iormac = io_iormac_213; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_214_clock = clock;
  assign bc_pe_214_reset = reset;
  assign bc_pe_214_io_ho_input = bc_pe_213_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_214_io_ve_input = bc_pe_198_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_214_io_input_valid = io_input_valid_214; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_214_io_iormac = io_iormac_214; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_215_clock = clock;
  assign bc_pe_215_reset = reset;
  assign bc_pe_215_io_ho_input = bc_pe_214_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_215_io_ve_input = bc_pe_199_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_215_io_input_valid = io_input_valid_215; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_215_io_iormac = io_iormac_215; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_216_clock = clock;
  assign bc_pe_216_reset = reset;
  assign bc_pe_216_io_ho_input = bc_pe_215_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_216_io_ve_input = bc_pe_200_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_216_io_input_valid = io_input_valid_216; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_216_io_iormac = io_iormac_216; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_217_clock = clock;
  assign bc_pe_217_reset = reset;
  assign bc_pe_217_io_ho_input = bc_pe_216_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_217_io_ve_input = bc_pe_201_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_217_io_input_valid = io_input_valid_217; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_217_io_iormac = io_iormac_217; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_218_clock = clock;
  assign bc_pe_218_reset = reset;
  assign bc_pe_218_io_ho_input = bc_pe_217_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_218_io_ve_input = bc_pe_202_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_218_io_input_valid = io_input_valid_218; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_218_io_iormac = io_iormac_218; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_219_clock = clock;
  assign bc_pe_219_reset = reset;
  assign bc_pe_219_io_ho_input = bc_pe_218_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_219_io_ve_input = bc_pe_203_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_219_io_input_valid = io_input_valid_219; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_219_io_iormac = io_iormac_219; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_220_clock = clock;
  assign bc_pe_220_reset = reset;
  assign bc_pe_220_io_ho_input = bc_pe_219_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_220_io_ve_input = bc_pe_204_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_220_io_input_valid = io_input_valid_220; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_220_io_iormac = io_iormac_220; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_221_clock = clock;
  assign bc_pe_221_reset = reset;
  assign bc_pe_221_io_ho_input = bc_pe_220_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_221_io_ve_input = bc_pe_205_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_221_io_input_valid = io_input_valid_221; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_221_io_iormac = io_iormac_221; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_222_clock = clock;
  assign bc_pe_222_reset = reset;
  assign bc_pe_222_io_ho_input = bc_pe_221_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_222_io_ve_input = bc_pe_206_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_222_io_input_valid = io_input_valid_222; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_222_io_iormac = io_iormac_222; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_223_clock = clock;
  assign bc_pe_223_reset = reset;
  assign bc_pe_223_io_ho_input = bc_pe_222_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_223_io_ve_input = bc_pe_207_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_223_io_input_valid = io_input_valid_223; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_223_io_iormac = io_iormac_223; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_224_clock = clock;
  assign bc_pe_224_reset = reset;
  assign bc_pe_224_io_ho_input = io_x_input_14; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_224_io_ve_input = bc_pe_208_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_224_io_input_valid = io_input_valid_224; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_224_io_iormac = io_iormac_224; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_225_clock = clock;
  assign bc_pe_225_reset = reset;
  assign bc_pe_225_io_ho_input = bc_pe_224_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_225_io_ve_input = bc_pe_209_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_225_io_input_valid = io_input_valid_225; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_225_io_iormac = io_iormac_225; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_226_clock = clock;
  assign bc_pe_226_reset = reset;
  assign bc_pe_226_io_ho_input = bc_pe_225_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_226_io_ve_input = bc_pe_210_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_226_io_input_valid = io_input_valid_226; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_226_io_iormac = io_iormac_226; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_227_clock = clock;
  assign bc_pe_227_reset = reset;
  assign bc_pe_227_io_ho_input = bc_pe_226_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_227_io_ve_input = bc_pe_211_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_227_io_input_valid = io_input_valid_227; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_227_io_iormac = io_iormac_227; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_228_clock = clock;
  assign bc_pe_228_reset = reset;
  assign bc_pe_228_io_ho_input = bc_pe_227_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_228_io_ve_input = bc_pe_212_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_228_io_input_valid = io_input_valid_228; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_228_io_iormac = io_iormac_228; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_229_clock = clock;
  assign bc_pe_229_reset = reset;
  assign bc_pe_229_io_ho_input = bc_pe_228_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_229_io_ve_input = bc_pe_213_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_229_io_input_valid = io_input_valid_229; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_229_io_iormac = io_iormac_229; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_230_clock = clock;
  assign bc_pe_230_reset = reset;
  assign bc_pe_230_io_ho_input = bc_pe_229_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_230_io_ve_input = bc_pe_214_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_230_io_input_valid = io_input_valid_230; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_230_io_iormac = io_iormac_230; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_231_clock = clock;
  assign bc_pe_231_reset = reset;
  assign bc_pe_231_io_ho_input = bc_pe_230_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_231_io_ve_input = bc_pe_215_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_231_io_input_valid = io_input_valid_231; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_231_io_iormac = io_iormac_231; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_232_clock = clock;
  assign bc_pe_232_reset = reset;
  assign bc_pe_232_io_ho_input = bc_pe_231_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_232_io_ve_input = bc_pe_216_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_232_io_input_valid = io_input_valid_232; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_232_io_iormac = io_iormac_232; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_233_clock = clock;
  assign bc_pe_233_reset = reset;
  assign bc_pe_233_io_ho_input = bc_pe_232_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_233_io_ve_input = bc_pe_217_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_233_io_input_valid = io_input_valid_233; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_233_io_iormac = io_iormac_233; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_234_clock = clock;
  assign bc_pe_234_reset = reset;
  assign bc_pe_234_io_ho_input = bc_pe_233_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_234_io_ve_input = bc_pe_218_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_234_io_input_valid = io_input_valid_234; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_234_io_iormac = io_iormac_234; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_235_clock = clock;
  assign bc_pe_235_reset = reset;
  assign bc_pe_235_io_ho_input = bc_pe_234_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_235_io_ve_input = bc_pe_219_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_235_io_input_valid = io_input_valid_235; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_235_io_iormac = io_iormac_235; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_236_clock = clock;
  assign bc_pe_236_reset = reset;
  assign bc_pe_236_io_ho_input = bc_pe_235_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_236_io_ve_input = bc_pe_220_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_236_io_input_valid = io_input_valid_236; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_236_io_iormac = io_iormac_236; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_237_clock = clock;
  assign bc_pe_237_reset = reset;
  assign bc_pe_237_io_ho_input = bc_pe_236_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_237_io_ve_input = bc_pe_221_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_237_io_input_valid = io_input_valid_237; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_237_io_iormac = io_iormac_237; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_238_clock = clock;
  assign bc_pe_238_reset = reset;
  assign bc_pe_238_io_ho_input = bc_pe_237_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_238_io_ve_input = bc_pe_222_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_238_io_input_valid = io_input_valid_238; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_238_io_iormac = io_iormac_238; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_239_clock = clock;
  assign bc_pe_239_reset = reset;
  assign bc_pe_239_io_ho_input = bc_pe_238_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_239_io_ve_input = bc_pe_223_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_239_io_input_valid = io_input_valid_239; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_239_io_iormac = io_iormac_239; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_240_clock = clock;
  assign bc_pe_240_reset = reset;
  assign bc_pe_240_io_ho_input = io_x_input_15; // @[bc_mmul.scala 22:28 60:41]
  assign bc_pe_240_io_ve_input = bc_pe_224_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_240_io_input_valid = io_input_valid_240; // @[bc_mmul.scala 22:28 62:41]
  assign bc_pe_240_io_iormac = io_iormac_240; // @[bc_mmul.scala 22:28 63:41]
  assign bc_pe_241_clock = clock;
  assign bc_pe_241_reset = reset;
  assign bc_pe_241_io_ho_input = bc_pe_240_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_241_io_ve_input = bc_pe_225_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_241_io_input_valid = io_input_valid_241; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_241_io_iormac = io_iormac_241; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_242_clock = clock;
  assign bc_pe_242_reset = reset;
  assign bc_pe_242_io_ho_input = bc_pe_241_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_242_io_ve_input = bc_pe_226_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_242_io_input_valid = io_input_valid_242; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_242_io_iormac = io_iormac_242; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_243_clock = clock;
  assign bc_pe_243_reset = reset;
  assign bc_pe_243_io_ho_input = bc_pe_242_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_243_io_ve_input = bc_pe_227_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_243_io_input_valid = io_input_valid_243; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_243_io_iormac = io_iormac_243; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_244_clock = clock;
  assign bc_pe_244_reset = reset;
  assign bc_pe_244_io_ho_input = bc_pe_243_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_244_io_ve_input = bc_pe_228_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_244_io_input_valid = io_input_valid_244; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_244_io_iormac = io_iormac_244; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_245_clock = clock;
  assign bc_pe_245_reset = reset;
  assign bc_pe_245_io_ho_input = bc_pe_244_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_245_io_ve_input = bc_pe_229_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_245_io_input_valid = io_input_valid_245; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_245_io_iormac = io_iormac_245; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_246_clock = clock;
  assign bc_pe_246_reset = reset;
  assign bc_pe_246_io_ho_input = bc_pe_245_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_246_io_ve_input = bc_pe_230_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_246_io_input_valid = io_input_valid_246; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_246_io_iormac = io_iormac_246; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_247_clock = clock;
  assign bc_pe_247_reset = reset;
  assign bc_pe_247_io_ho_input = bc_pe_246_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_247_io_ve_input = bc_pe_231_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_247_io_input_valid = io_input_valid_247; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_247_io_iormac = io_iormac_247; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_248_clock = clock;
  assign bc_pe_248_reset = reset;
  assign bc_pe_248_io_ho_input = bc_pe_247_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_248_io_ve_input = bc_pe_232_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_248_io_input_valid = io_input_valid_248; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_248_io_iormac = io_iormac_248; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_249_clock = clock;
  assign bc_pe_249_reset = reset;
  assign bc_pe_249_io_ho_input = bc_pe_248_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_249_io_ve_input = bc_pe_233_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_249_io_input_valid = io_input_valid_249; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_249_io_iormac = io_iormac_249; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_250_clock = clock;
  assign bc_pe_250_reset = reset;
  assign bc_pe_250_io_ho_input = bc_pe_249_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_250_io_ve_input = bc_pe_234_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_250_io_input_valid = io_input_valid_250; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_250_io_iormac = io_iormac_250; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_251_clock = clock;
  assign bc_pe_251_reset = reset;
  assign bc_pe_251_io_ho_input = bc_pe_250_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_251_io_ve_input = bc_pe_235_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_251_io_input_valid = io_input_valid_251; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_251_io_iormac = io_iormac_251; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_252_clock = clock;
  assign bc_pe_252_reset = reset;
  assign bc_pe_252_io_ho_input = bc_pe_251_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_252_io_ve_input = bc_pe_236_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_252_io_input_valid = io_input_valid_252; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_252_io_iormac = io_iormac_252; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_253_clock = clock;
  assign bc_pe_253_reset = reset;
  assign bc_pe_253_io_ho_input = bc_pe_252_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_253_io_ve_input = bc_pe_237_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_253_io_input_valid = io_input_valid_253; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_253_io_iormac = io_iormac_253; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_254_clock = clock;
  assign bc_pe_254_reset = reset;
  assign bc_pe_254_io_ho_input = bc_pe_253_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_254_io_ve_input = bc_pe_238_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_254_io_input_valid = io_input_valid_254; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_254_io_iormac = io_iormac_254; // @[bc_mmul.scala 22:28 78:47]
  assign bc_pe_255_clock = clock;
  assign bc_pe_255_reset = reset;
  assign bc_pe_255_io_ho_input = bc_pe_254_io_ho_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_255_io_ve_input = bc_pe_239_io_ve_out; // @[bc_mmul.scala 22:{28,28}]
  assign bc_pe_255_io_input_valid = io_input_valid_255; // @[bc_mmul.scala 22:28 77:47]
  assign bc_pe_255_io_iormac = io_iormac_255; // @[bc_mmul.scala 22:28 78:47]
endmodule
